module magic_mem
(
	input logic clk,
	input logic reset,
	
	// Row select
	input logic [31:0] row_sel,
	
	// Output row
	output logic [31:0] row[63:0]
);

	logic [31:0] data[63:0][63:0]; // 64x64 FP array
	logic [31:0] row_reg[63:0];    // Holds selected row
	
	// Assign 64 * i + j
	initial begin
        data[0][0] = 32'h0;
        data[0][1] = 32'h3f800000;
        data[0][2] = 32'h40000000;
        data[0][3] = 32'h40400000;
        data[0][4] = 32'h40800000;
        data[0][5] = 32'h40a00000;
        data[0][6] = 32'h40c00000;
        data[0][7] = 32'h40e00000;
        data[0][8] = 32'h41000000;
        data[0][9] = 32'h41100000;
        data[0][10] = 32'h41200000;
        data[0][11] = 32'h41300000;
        data[0][12] = 32'h41400000;
        data[0][13] = 32'h41500000;
        data[0][14] = 32'h41600000;
        data[0][15] = 32'h41700000;
        data[0][16] = 32'h41800000;
        data[0][17] = 32'h41880000;
        data[0][18] = 32'h41900000;
        data[0][19] = 32'h41980000;
        data[0][20] = 32'h41a00000;
        data[0][21] = 32'h41a80000;
        data[0][22] = 32'h41b00000;
        data[0][23] = 32'h41b80000;
        data[0][24] = 32'h41c00000;
        data[0][25] = 32'h41c80000;
        data[0][26] = 32'h41d00000;
        data[0][27] = 32'h41d80000;
        data[0][28] = 32'h41e00000;
        data[0][29] = 32'h41e80000;
        data[0][30] = 32'h41f00000;
        data[0][31] = 32'h41f80000;
        data[0][32] = 32'h42000000;
        data[0][33] = 32'h42040000;
        data[0][34] = 32'h42080000;
        data[0][35] = 32'h420c0000;
        data[0][36] = 32'h42100000;
        data[0][37] = 32'h42140000;
        data[0][38] = 32'h42180000;
        data[0][39] = 32'h421c0000;
        data[0][40] = 32'h42200000;
        data[0][41] = 32'h42240000;
        data[0][42] = 32'h42280000;
        data[0][43] = 32'h422c0000;
        data[0][44] = 32'h42300000;
        data[0][45] = 32'h42340000;
        data[0][46] = 32'h42380000;
        data[0][47] = 32'h423c0000;
        data[0][48] = 32'h42400000;
        data[0][49] = 32'h42440000;
        data[0][50] = 32'h42480000;
        data[0][51] = 32'h424c0000;
        data[0][52] = 32'h42500000;
        data[0][53] = 32'h42540000;
        data[0][54] = 32'h42580000;
        data[0][55] = 32'h425c0000;
        data[0][56] = 32'h42600000;
        data[0][57] = 32'h42640000;
        data[0][58] = 32'h42680000;
        data[0][59] = 32'h426c0000;
        data[0][60] = 32'h42700000;
        data[0][61] = 32'h42740000;
        data[0][62] = 32'h42780000;
        data[0][63] = 32'h427c0000;
        data[1][0] = 32'h42800000;
        data[1][1] = 32'h42820000;
        data[1][2] = 32'h42840000;
        data[1][3] = 32'h42860000;
        data[1][4] = 32'h42880000;
        data[1][5] = 32'h428a0000;
        data[1][6] = 32'h428c0000;
        data[1][7] = 32'h428e0000;
        data[1][8] = 32'h42900000;
        data[1][9] = 32'h42920000;
        data[1][10] = 32'h42940000;
        data[1][11] = 32'h42960000;
        data[1][12] = 32'h42980000;
        data[1][13] = 32'h429a0000;
        data[1][14] = 32'h429c0000;
        data[1][15] = 32'h429e0000;
        data[1][16] = 32'h42a00000;
        data[1][17] = 32'h42a20000;
        data[1][18] = 32'h42a40000;
        data[1][19] = 32'h42a60000;
        data[1][20] = 32'h42a80000;
        data[1][21] = 32'h42aa0000;
        data[1][22] = 32'h42ac0000;
        data[1][23] = 32'h42ae0000;
        data[1][24] = 32'h42b00000;
        data[1][25] = 32'h42b20000;
        data[1][26] = 32'h42b40000;
        data[1][27] = 32'h42b60000;
        data[1][28] = 32'h42b80000;
        data[1][29] = 32'h42ba0000;
        data[1][30] = 32'h42bc0000;
        data[1][31] = 32'h42be0000;
        data[1][32] = 32'h42c00000;
        data[1][33] = 32'h42c20000;
        data[1][34] = 32'h42c40000;
        data[1][35] = 32'h42c60000;
        data[1][36] = 32'h42c80000;
        data[1][37] = 32'h42ca0000;
        data[1][38] = 32'h42cc0000;
        data[1][39] = 32'h42ce0000;
        data[1][40] = 32'h42d00000;
        data[1][41] = 32'h42d20000;
        data[1][42] = 32'h42d40000;
        data[1][43] = 32'h42d60000;
        data[1][44] = 32'h42d80000;
        data[1][45] = 32'h42da0000;
        data[1][46] = 32'h42dc0000;
        data[1][47] = 32'h42de0000;
        data[1][48] = 32'h42e00000;
        data[1][49] = 32'h42e20000;
        data[1][50] = 32'h42e40000;
        data[1][51] = 32'h42e60000;
        data[1][52] = 32'h42e80000;
        data[1][53] = 32'h42ea0000;
        data[1][54] = 32'h42ec0000;
        data[1][55] = 32'h42ee0000;
        data[1][56] = 32'h42f00000;
        data[1][57] = 32'h42f20000;
        data[1][58] = 32'h42f40000;
        data[1][59] = 32'h42f60000;
        data[1][60] = 32'h42f80000;
        data[1][61] = 32'h42fa0000;
        data[1][62] = 32'h42fc0000;
        data[1][63] = 32'h42fe0000;
        data[2][0] = 32'h43000000;
        data[2][1] = 32'h43010000;
        data[2][2] = 32'h43020000;
        data[2][3] = 32'h43030000;
        data[2][4] = 32'h43040000;
        data[2][5] = 32'h43050000;
        data[2][6] = 32'h43060000;
        data[2][7] = 32'h43070000;
        data[2][8] = 32'h43080000;
        data[2][9] = 32'h43090000;
        data[2][10] = 32'h430a0000;
        data[2][11] = 32'h430b0000;
        data[2][12] = 32'h430c0000;
        data[2][13] = 32'h430d0000;
        data[2][14] = 32'h430e0000;
        data[2][15] = 32'h430f0000;
        data[2][16] = 32'h43100000;
        data[2][17] = 32'h43110000;
        data[2][18] = 32'h43120000;
        data[2][19] = 32'h43130000;
        data[2][20] = 32'h43140000;
        data[2][21] = 32'h43150000;
        data[2][22] = 32'h43160000;
        data[2][23] = 32'h43170000;
        data[2][24] = 32'h43180000;
        data[2][25] = 32'h43190000;
        data[2][26] = 32'h431a0000;
        data[2][27] = 32'h431b0000;
        data[2][28] = 32'h431c0000;
        data[2][29] = 32'h431d0000;
        data[2][30] = 32'h431e0000;
        data[2][31] = 32'h431f0000;
        data[2][32] = 32'h43200000;
        data[2][33] = 32'h43210000;
        data[2][34] = 32'h43220000;
        data[2][35] = 32'h43230000;
        data[2][36] = 32'h43240000;
        data[2][37] = 32'h43250000;
        data[2][38] = 32'h43260000;
        data[2][39] = 32'h43270000;
        data[2][40] = 32'h43280000;
        data[2][41] = 32'h43290000;
        data[2][42] = 32'h432a0000;
        data[2][43] = 32'h432b0000;
        data[2][44] = 32'h432c0000;
        data[2][45] = 32'h432d0000;
        data[2][46] = 32'h432e0000;
        data[2][47] = 32'h432f0000;
        data[2][48] = 32'h43300000;
        data[2][49] = 32'h43310000;
        data[2][50] = 32'h43320000;
        data[2][51] = 32'h43330000;
        data[2][52] = 32'h43340000;
        data[2][53] = 32'h43350000;
        data[2][54] = 32'h43360000;
        data[2][55] = 32'h43370000;
        data[2][56] = 32'h43380000;
        data[2][57] = 32'h43390000;
        data[2][58] = 32'h433a0000;
        data[2][59] = 32'h433b0000;
        data[2][60] = 32'h433c0000;
        data[2][61] = 32'h433d0000;
        data[2][62] = 32'h433e0000;
        data[2][63] = 32'h433f0000;
        data[3][0] = 32'h43400000;
        data[3][1] = 32'h43410000;
        data[3][2] = 32'h43420000;
        data[3][3] = 32'h43430000;
        data[3][4] = 32'h43440000;
        data[3][5] = 32'h43450000;
        data[3][6] = 32'h43460000;
        data[3][7] = 32'h43470000;
        data[3][8] = 32'h43480000;
        data[3][9] = 32'h43490000;
        data[3][10] = 32'h434a0000;
        data[3][11] = 32'h434b0000;
        data[3][12] = 32'h434c0000;
        data[3][13] = 32'h434d0000;
        data[3][14] = 32'h434e0000;
        data[3][15] = 32'h434f0000;
        data[3][16] = 32'h43500000;
        data[3][17] = 32'h43510000;
        data[3][18] = 32'h43520000;
        data[3][19] = 32'h43530000;
        data[3][20] = 32'h43540000;
        data[3][21] = 32'h43550000;
        data[3][22] = 32'h43560000;
        data[3][23] = 32'h43570000;
        data[3][24] = 32'h43580000;
        data[3][25] = 32'h43590000;
        data[3][26] = 32'h435a0000;
        data[3][27] = 32'h435b0000;
        data[3][28] = 32'h435c0000;
        data[3][29] = 32'h435d0000;
        data[3][30] = 32'h435e0000;
        data[3][31] = 32'h435f0000;
        data[3][32] = 32'h43600000;
        data[3][33] = 32'h43610000;
        data[3][34] = 32'h43620000;
        data[3][35] = 32'h43630000;
        data[3][36] = 32'h43640000;
        data[3][37] = 32'h43650000;
        data[3][38] = 32'h43660000;
        data[3][39] = 32'h43670000;
        data[3][40] = 32'h43680000;
        data[3][41] = 32'h43690000;
        data[3][42] = 32'h436a0000;
        data[3][43] = 32'h436b0000;
        data[3][44] = 32'h436c0000;
        data[3][45] = 32'h436d0000;
        data[3][46] = 32'h436e0000;
        data[3][47] = 32'h436f0000;
        data[3][48] = 32'h43700000;
        data[3][49] = 32'h43710000;
        data[3][50] = 32'h43720000;
        data[3][51] = 32'h43730000;
        data[3][52] = 32'h43740000;
        data[3][53] = 32'h43750000;
        data[3][54] = 32'h43760000;
        data[3][55] = 32'h43770000;
        data[3][56] = 32'h43780000;
        data[3][57] = 32'h43790000;
        data[3][58] = 32'h437a0000;
        data[3][59] = 32'h437b0000;
        data[3][60] = 32'h437c0000;
        data[3][61] = 32'h437d0000;
        data[3][62] = 32'h437e0000;
        data[3][63] = 32'h437f0000;
        data[4][0] = 32'h43800000;
        data[4][1] = 32'h43808000;
        data[4][2] = 32'h43810000;
        data[4][3] = 32'h43818000;
        data[4][4] = 32'h43820000;
        data[4][5] = 32'h43828000;
        data[4][6] = 32'h43830000;
        data[4][7] = 32'h43838000;
        data[4][8] = 32'h43840000;
        data[4][9] = 32'h43848000;
        data[4][10] = 32'h43850000;
        data[4][11] = 32'h43858000;
        data[4][12] = 32'h43860000;
        data[4][13] = 32'h43868000;
        data[4][14] = 32'h43870000;
        data[4][15] = 32'h43878000;
        data[4][16] = 32'h43880000;
        data[4][17] = 32'h43888000;
        data[4][18] = 32'h43890000;
        data[4][19] = 32'h43898000;
        data[4][20] = 32'h438a0000;
        data[4][21] = 32'h438a8000;
        data[4][22] = 32'h438b0000;
        data[4][23] = 32'h438b8000;
        data[4][24] = 32'h438c0000;
        data[4][25] = 32'h438c8000;
        data[4][26] = 32'h438d0000;
        data[4][27] = 32'h438d8000;
        data[4][28] = 32'h438e0000;
        data[4][29] = 32'h438e8000;
        data[4][30] = 32'h438f0000;
        data[4][31] = 32'h438f8000;
        data[4][32] = 32'h43900000;
        data[4][33] = 32'h43908000;
        data[4][34] = 32'h43910000;
        data[4][35] = 32'h43918000;
        data[4][36] = 32'h43920000;
        data[4][37] = 32'h43928000;
        data[4][38] = 32'h43930000;
        data[4][39] = 32'h43938000;
        data[4][40] = 32'h43940000;
        data[4][41] = 32'h43948000;
        data[4][42] = 32'h43950000;
        data[4][43] = 32'h43958000;
        data[4][44] = 32'h43960000;
        data[4][45] = 32'h43968000;
        data[4][46] = 32'h43970000;
        data[4][47] = 32'h43978000;
        data[4][48] = 32'h43980000;
        data[4][49] = 32'h43988000;
        data[4][50] = 32'h43990000;
        data[4][51] = 32'h43998000;
        data[4][52] = 32'h439a0000;
        data[4][53] = 32'h439a8000;
        data[4][54] = 32'h439b0000;
        data[4][55] = 32'h439b8000;
        data[4][56] = 32'h439c0000;
        data[4][57] = 32'h439c8000;
        data[4][58] = 32'h439d0000;
        data[4][59] = 32'h439d8000;
        data[4][60] = 32'h439e0000;
        data[4][61] = 32'h439e8000;
        data[4][62] = 32'h439f0000;
        data[4][63] = 32'h439f8000;
        data[5][0] = 32'h43a00000;
        data[5][1] = 32'h43a08000;
        data[5][2] = 32'h43a10000;
        data[5][3] = 32'h43a18000;
        data[5][4] = 32'h43a20000;
        data[5][5] = 32'h43a28000;
        data[5][6] = 32'h43a30000;
        data[5][7] = 32'h43a38000;
        data[5][8] = 32'h43a40000;
        data[5][9] = 32'h43a48000;
        data[5][10] = 32'h43a50000;
        data[5][11] = 32'h43a58000;
        data[5][12] = 32'h43a60000;
        data[5][13] = 32'h43a68000;
        data[5][14] = 32'h43a70000;
        data[5][15] = 32'h43a78000;
        data[5][16] = 32'h43a80000;
        data[5][17] = 32'h43a88000;
        data[5][18] = 32'h43a90000;
        data[5][19] = 32'h43a98000;
        data[5][20] = 32'h43aa0000;
        data[5][21] = 32'h43aa8000;
        data[5][22] = 32'h43ab0000;
        data[5][23] = 32'h43ab8000;
        data[5][24] = 32'h43ac0000;
        data[5][25] = 32'h43ac8000;
        data[5][26] = 32'h43ad0000;
        data[5][27] = 32'h43ad8000;
        data[5][28] = 32'h43ae0000;
        data[5][29] = 32'h43ae8000;
        data[5][30] = 32'h43af0000;
        data[5][31] = 32'h43af8000;
        data[5][32] = 32'h43b00000;
        data[5][33] = 32'h43b08000;
        data[5][34] = 32'h43b10000;
        data[5][35] = 32'h43b18000;
        data[5][36] = 32'h43b20000;
        data[5][37] = 32'h43b28000;
        data[5][38] = 32'h43b30000;
        data[5][39] = 32'h43b38000;
        data[5][40] = 32'h43b40000;
        data[5][41] = 32'h43b48000;
        data[5][42] = 32'h43b50000;
        data[5][43] = 32'h43b58000;
        data[5][44] = 32'h43b60000;
        data[5][45] = 32'h43b68000;
        data[5][46] = 32'h43b70000;
        data[5][47] = 32'h43b78000;
        data[5][48] = 32'h43b80000;
        data[5][49] = 32'h43b88000;
        data[5][50] = 32'h43b90000;
        data[5][51] = 32'h43b98000;
        data[5][52] = 32'h43ba0000;
        data[5][53] = 32'h43ba8000;
        data[5][54] = 32'h43bb0000;
        data[5][55] = 32'h43bb8000;
        data[5][56] = 32'h43bc0000;
        data[5][57] = 32'h43bc8000;
        data[5][58] = 32'h43bd0000;
        data[5][59] = 32'h43bd8000;
        data[5][60] = 32'h43be0000;
        data[5][61] = 32'h43be8000;
        data[5][62] = 32'h43bf0000;
        data[5][63] = 32'h43bf8000;
        data[6][0] = 32'h43c00000;
        data[6][1] = 32'h43c08000;
        data[6][2] = 32'h43c10000;
        data[6][3] = 32'h43c18000;
        data[6][4] = 32'h43c20000;
        data[6][5] = 32'h43c28000;
        data[6][6] = 32'h43c30000;
        data[6][7] = 32'h43c38000;
        data[6][8] = 32'h43c40000;
        data[6][9] = 32'h43c48000;
        data[6][10] = 32'h43c50000;
        data[6][11] = 32'h43c58000;
        data[6][12] = 32'h43c60000;
        data[6][13] = 32'h43c68000;
        data[6][14] = 32'h43c70000;
        data[6][15] = 32'h43c78000;
        data[6][16] = 32'h43c80000;
        data[6][17] = 32'h43c88000;
        data[6][18] = 32'h43c90000;
        data[6][19] = 32'h43c98000;
        data[6][20] = 32'h43ca0000;
        data[6][21] = 32'h43ca8000;
        data[6][22] = 32'h43cb0000;
        data[6][23] = 32'h43cb8000;
        data[6][24] = 32'h43cc0000;
        data[6][25] = 32'h43cc8000;
        data[6][26] = 32'h43cd0000;
        data[6][27] = 32'h43cd8000;
        data[6][28] = 32'h43ce0000;
        data[6][29] = 32'h43ce8000;
        data[6][30] = 32'h43cf0000;
        data[6][31] = 32'h43cf8000;
        data[6][32] = 32'h43d00000;
        data[6][33] = 32'h43d08000;
        data[6][34] = 32'h43d10000;
        data[6][35] = 32'h43d18000;
        data[6][36] = 32'h43d20000;
        data[6][37] = 32'h43d28000;
        data[6][38] = 32'h43d30000;
        data[6][39] = 32'h43d38000;
        data[6][40] = 32'h43d40000;
        data[6][41] = 32'h43d48000;
        data[6][42] = 32'h43d50000;
        data[6][43] = 32'h43d58000;
        data[6][44] = 32'h43d60000;
        data[6][45] = 32'h43d68000;
        data[6][46] = 32'h43d70000;
        data[6][47] = 32'h43d78000;
        data[6][48] = 32'h43d80000;
        data[6][49] = 32'h43d88000;
        data[6][50] = 32'h43d90000;
        data[6][51] = 32'h43d98000;
        data[6][52] = 32'h43da0000;
        data[6][53] = 32'h43da8000;
        data[6][54] = 32'h43db0000;
        data[6][55] = 32'h43db8000;
        data[6][56] = 32'h43dc0000;
        data[6][57] = 32'h43dc8000;
        data[6][58] = 32'h43dd0000;
        data[6][59] = 32'h43dd8000;
        data[6][60] = 32'h43de0000;
        data[6][61] = 32'h43de8000;
        data[6][62] = 32'h43df0000;
        data[6][63] = 32'h43df8000;
        data[7][0] = 32'h43e00000;
        data[7][1] = 32'h43e08000;
        data[7][2] = 32'h43e10000;
        data[7][3] = 32'h43e18000;
        data[7][4] = 32'h43e20000;
        data[7][5] = 32'h43e28000;
        data[7][6] = 32'h43e30000;
        data[7][7] = 32'h43e38000;
        data[7][8] = 32'h43e40000;
        data[7][9] = 32'h43e48000;
        data[7][10] = 32'h43e50000;
        data[7][11] = 32'h43e58000;
        data[7][12] = 32'h43e60000;
        data[7][13] = 32'h43e68000;
        data[7][14] = 32'h43e70000;
        data[7][15] = 32'h43e78000;
        data[7][16] = 32'h43e80000;
        data[7][17] = 32'h43e88000;
        data[7][18] = 32'h43e90000;
        data[7][19] = 32'h43e98000;
        data[7][20] = 32'h43ea0000;
        data[7][21] = 32'h43ea8000;
        data[7][22] = 32'h43eb0000;
        data[7][23] = 32'h43eb8000;
        data[7][24] = 32'h43ec0000;
        data[7][25] = 32'h43ec8000;
        data[7][26] = 32'h43ed0000;
        data[7][27] = 32'h43ed8000;
        data[7][28] = 32'h43ee0000;
        data[7][29] = 32'h43ee8000;
        data[7][30] = 32'h43ef0000;
        data[7][31] = 32'h43ef8000;
        data[7][32] = 32'h43f00000;
        data[7][33] = 32'h43f08000;
        data[7][34] = 32'h43f10000;
        data[7][35] = 32'h43f18000;
        data[7][36] = 32'h43f20000;
        data[7][37] = 32'h43f28000;
        data[7][38] = 32'h43f30000;
        data[7][39] = 32'h43f38000;
        data[7][40] = 32'h43f40000;
        data[7][41] = 32'h43f48000;
        data[7][42] = 32'h43f50000;
        data[7][43] = 32'h43f58000;
        data[7][44] = 32'h43f60000;
        data[7][45] = 32'h43f68000;
        data[7][46] = 32'h43f70000;
        data[7][47] = 32'h43f78000;
        data[7][48] = 32'h43f80000;
        data[7][49] = 32'h43f88000;
        data[7][50] = 32'h43f90000;
        data[7][51] = 32'h43f98000;
        data[7][52] = 32'h43fa0000;
        data[7][53] = 32'h43fa8000;
        data[7][54] = 32'h43fb0000;
        data[7][55] = 32'h43fb8000;
        data[7][56] = 32'h43fc0000;
        data[7][57] = 32'h43fc8000;
        data[7][58] = 32'h43fd0000;
        data[7][59] = 32'h43fd8000;
        data[7][60] = 32'h43fe0000;
        data[7][61] = 32'h43fe8000;
        data[7][62] = 32'h43ff0000;
        data[7][63] = 32'h43ff8000;
        data[8][0] = 32'h44000000;
        data[8][1] = 32'h44004000;
        data[8][2] = 32'h44008000;
        data[8][3] = 32'h4400c000;
        data[8][4] = 32'h44010000;
        data[8][5] = 32'h44014000;
        data[8][6] = 32'h44018000;
        data[8][7] = 32'h4401c000;
        data[8][8] = 32'h44020000;
        data[8][9] = 32'h44024000;
        data[8][10] = 32'h44028000;
        data[8][11] = 32'h4402c000;
        data[8][12] = 32'h44030000;
        data[8][13] = 32'h44034000;
        data[8][14] = 32'h44038000;
        data[8][15] = 32'h4403c000;
        data[8][16] = 32'h44040000;
        data[8][17] = 32'h44044000;
        data[8][18] = 32'h44048000;
        data[8][19] = 32'h4404c000;
        data[8][20] = 32'h44050000;
        data[8][21] = 32'h44054000;
        data[8][22] = 32'h44058000;
        data[8][23] = 32'h4405c000;
        data[8][24] = 32'h44060000;
        data[8][25] = 32'h44064000;
        data[8][26] = 32'h44068000;
        data[8][27] = 32'h4406c000;
        data[8][28] = 32'h44070000;
        data[8][29] = 32'h44074000;
        data[8][30] = 32'h44078000;
        data[8][31] = 32'h4407c000;
        data[8][32] = 32'h44080000;
        data[8][33] = 32'h44084000;
        data[8][34] = 32'h44088000;
        data[8][35] = 32'h4408c000;
        data[8][36] = 32'h44090000;
        data[8][37] = 32'h44094000;
        data[8][38] = 32'h44098000;
        data[8][39] = 32'h4409c000;
        data[8][40] = 32'h440a0000;
        data[8][41] = 32'h440a4000;
        data[8][42] = 32'h440a8000;
        data[8][43] = 32'h440ac000;
        data[8][44] = 32'h440b0000;
        data[8][45] = 32'h440b4000;
        data[8][46] = 32'h440b8000;
        data[8][47] = 32'h440bc000;
        data[8][48] = 32'h440c0000;
        data[8][49] = 32'h440c4000;
        data[8][50] = 32'h440c8000;
        data[8][51] = 32'h440cc000;
        data[8][52] = 32'h440d0000;
        data[8][53] = 32'h440d4000;
        data[8][54] = 32'h440d8000;
        data[8][55] = 32'h440dc000;
        data[8][56] = 32'h440e0000;
        data[8][57] = 32'h440e4000;
        data[8][58] = 32'h440e8000;
        data[8][59] = 32'h440ec000;
        data[8][60] = 32'h440f0000;
        data[8][61] = 32'h440f4000;
        data[8][62] = 32'h440f8000;
        data[8][63] = 32'h440fc000;
        data[9][0] = 32'h44100000;
        data[9][1] = 32'h44104000;
        data[9][2] = 32'h44108000;
        data[9][3] = 32'h4410c000;
        data[9][4] = 32'h44110000;
        data[9][5] = 32'h44114000;
        data[9][6] = 32'h44118000;
        data[9][7] = 32'h4411c000;
        data[9][8] = 32'h44120000;
        data[9][9] = 32'h44124000;
        data[9][10] = 32'h44128000;
        data[9][11] = 32'h4412c000;
        data[9][12] = 32'h44130000;
        data[9][13] = 32'h44134000;
        data[9][14] = 32'h44138000;
        data[9][15] = 32'h4413c000;
        data[9][16] = 32'h44140000;
        data[9][17] = 32'h44144000;
        data[9][18] = 32'h44148000;
        data[9][19] = 32'h4414c000;
        data[9][20] = 32'h44150000;
        data[9][21] = 32'h44154000;
        data[9][22] = 32'h44158000;
        data[9][23] = 32'h4415c000;
        data[9][24] = 32'h44160000;
        data[9][25] = 32'h44164000;
        data[9][26] = 32'h44168000;
        data[9][27] = 32'h4416c000;
        data[9][28] = 32'h44170000;
        data[9][29] = 32'h44174000;
        data[9][30] = 32'h44178000;
        data[9][31] = 32'h4417c000;
        data[9][32] = 32'h44180000;
        data[9][33] = 32'h44184000;
        data[9][34] = 32'h44188000;
        data[9][35] = 32'h4418c000;
        data[9][36] = 32'h44190000;
        data[9][37] = 32'h44194000;
        data[9][38] = 32'h44198000;
        data[9][39] = 32'h4419c000;
        data[9][40] = 32'h441a0000;
        data[9][41] = 32'h441a4000;
        data[9][42] = 32'h441a8000;
        data[9][43] = 32'h441ac000;
        data[9][44] = 32'h441b0000;
        data[9][45] = 32'h441b4000;
        data[9][46] = 32'h441b8000;
        data[9][47] = 32'h441bc000;
        data[9][48] = 32'h441c0000;
        data[9][49] = 32'h441c4000;
        data[9][50] = 32'h441c8000;
        data[9][51] = 32'h441cc000;
        data[9][52] = 32'h441d0000;
        data[9][53] = 32'h441d4000;
        data[9][54] = 32'h441d8000;
        data[9][55] = 32'h441dc000;
        data[9][56] = 32'h441e0000;
        data[9][57] = 32'h441e4000;
        data[9][58] = 32'h441e8000;
        data[9][59] = 32'h441ec000;
        data[9][60] = 32'h441f0000;
        data[9][61] = 32'h441f4000;
        data[9][62] = 32'h441f8000;
        data[9][63] = 32'h441fc000;
        data[10][0] = 32'h44200000;
        data[10][1] = 32'h44204000;
        data[10][2] = 32'h44208000;
        data[10][3] = 32'h4420c000;
        data[10][4] = 32'h44210000;
        data[10][5] = 32'h44214000;
        data[10][6] = 32'h44218000;
        data[10][7] = 32'h4421c000;
        data[10][8] = 32'h44220000;
        data[10][9] = 32'h44224000;
        data[10][10] = 32'h44228000;
        data[10][11] = 32'h4422c000;
        data[10][12] = 32'h44230000;
        data[10][13] = 32'h44234000;
        data[10][14] = 32'h44238000;
        data[10][15] = 32'h4423c000;
        data[10][16] = 32'h44240000;
        data[10][17] = 32'h44244000;
        data[10][18] = 32'h44248000;
        data[10][19] = 32'h4424c000;
        data[10][20] = 32'h44250000;
        data[10][21] = 32'h44254000;
        data[10][22] = 32'h44258000;
        data[10][23] = 32'h4425c000;
        data[10][24] = 32'h44260000;
        data[10][25] = 32'h44264000;
        data[10][26] = 32'h44268000;
        data[10][27] = 32'h4426c000;
        data[10][28] = 32'h44270000;
        data[10][29] = 32'h44274000;
        data[10][30] = 32'h44278000;
        data[10][31] = 32'h4427c000;
        data[10][32] = 32'h44280000;
        data[10][33] = 32'h44284000;
        data[10][34] = 32'h44288000;
        data[10][35] = 32'h4428c000;
        data[10][36] = 32'h44290000;
        data[10][37] = 32'h44294000;
        data[10][38] = 32'h44298000;
        data[10][39] = 32'h4429c000;
        data[10][40] = 32'h442a0000;
        data[10][41] = 32'h442a4000;
        data[10][42] = 32'h442a8000;
        data[10][43] = 32'h442ac000;
        data[10][44] = 32'h442b0000;
        data[10][45] = 32'h442b4000;
        data[10][46] = 32'h442b8000;
        data[10][47] = 32'h442bc000;
        data[10][48] = 32'h442c0000;
        data[10][49] = 32'h442c4000;
        data[10][50] = 32'h442c8000;
        data[10][51] = 32'h442cc000;
        data[10][52] = 32'h442d0000;
        data[10][53] = 32'h442d4000;
        data[10][54] = 32'h442d8000;
        data[10][55] = 32'h442dc000;
        data[10][56] = 32'h442e0000;
        data[10][57] = 32'h442e4000;
        data[10][58] = 32'h442e8000;
        data[10][59] = 32'h442ec000;
        data[10][60] = 32'h442f0000;
        data[10][61] = 32'h442f4000;
        data[10][62] = 32'h442f8000;
        data[10][63] = 32'h442fc000;
        data[11][0] = 32'h44300000;
        data[11][1] = 32'h44304000;
        data[11][2] = 32'h44308000;
        data[11][3] = 32'h4430c000;
        data[11][4] = 32'h44310000;
        data[11][5] = 32'h44314000;
        data[11][6] = 32'h44318000;
        data[11][7] = 32'h4431c000;
        data[11][8] = 32'h44320000;
        data[11][9] = 32'h44324000;
        data[11][10] = 32'h44328000;
        data[11][11] = 32'h4432c000;
        data[11][12] = 32'h44330000;
        data[11][13] = 32'h44334000;
        data[11][14] = 32'h44338000;
        data[11][15] = 32'h4433c000;
        data[11][16] = 32'h44340000;
        data[11][17] = 32'h44344000;
        data[11][18] = 32'h44348000;
        data[11][19] = 32'h4434c000;
        data[11][20] = 32'h44350000;
        data[11][21] = 32'h44354000;
        data[11][22] = 32'h44358000;
        data[11][23] = 32'h4435c000;
        data[11][24] = 32'h44360000;
        data[11][25] = 32'h44364000;
        data[11][26] = 32'h44368000;
        data[11][27] = 32'h4436c000;
        data[11][28] = 32'h44370000;
        data[11][29] = 32'h44374000;
        data[11][30] = 32'h44378000;
        data[11][31] = 32'h4437c000;
        data[11][32] = 32'h44380000;
        data[11][33] = 32'h44384000;
        data[11][34] = 32'h44388000;
        data[11][35] = 32'h4438c000;
        data[11][36] = 32'h44390000;
        data[11][37] = 32'h44394000;
        data[11][38] = 32'h44398000;
        data[11][39] = 32'h4439c000;
        data[11][40] = 32'h443a0000;
        data[11][41] = 32'h443a4000;
        data[11][42] = 32'h443a8000;
        data[11][43] = 32'h443ac000;
        data[11][44] = 32'h443b0000;
        data[11][45] = 32'h443b4000;
        data[11][46] = 32'h443b8000;
        data[11][47] = 32'h443bc000;
        data[11][48] = 32'h443c0000;
        data[11][49] = 32'h443c4000;
        data[11][50] = 32'h443c8000;
        data[11][51] = 32'h443cc000;
        data[11][52] = 32'h443d0000;
        data[11][53] = 32'h443d4000;
        data[11][54] = 32'h443d8000;
        data[11][55] = 32'h443dc000;
        data[11][56] = 32'h443e0000;
        data[11][57] = 32'h443e4000;
        data[11][58] = 32'h443e8000;
        data[11][59] = 32'h443ec000;
        data[11][60] = 32'h443f0000;
        data[11][61] = 32'h443f4000;
        data[11][62] = 32'h443f8000;
        data[11][63] = 32'h443fc000;
        data[12][0] = 32'h44400000;
        data[12][1] = 32'h44404000;
        data[12][2] = 32'h44408000;
        data[12][3] = 32'h4440c000;
        data[12][4] = 32'h44410000;
        data[12][5] = 32'h44414000;
        data[12][6] = 32'h44418000;
        data[12][7] = 32'h4441c000;
        data[12][8] = 32'h44420000;
        data[12][9] = 32'h44424000;
        data[12][10] = 32'h44428000;
        data[12][11] = 32'h4442c000;
        data[12][12] = 32'h44430000;
        data[12][13] = 32'h44434000;
        data[12][14] = 32'h44438000;
        data[12][15] = 32'h4443c000;
        data[12][16] = 32'h44440000;
        data[12][17] = 32'h44444000;
        data[12][18] = 32'h44448000;
        data[12][19] = 32'h4444c000;
        data[12][20] = 32'h44450000;
        data[12][21] = 32'h44454000;
        data[12][22] = 32'h44458000;
        data[12][23] = 32'h4445c000;
        data[12][24] = 32'h44460000;
        data[12][25] = 32'h44464000;
        data[12][26] = 32'h44468000;
        data[12][27] = 32'h4446c000;
        data[12][28] = 32'h44470000;
        data[12][29] = 32'h44474000;
        data[12][30] = 32'h44478000;
        data[12][31] = 32'h4447c000;
        data[12][32] = 32'h44480000;
        data[12][33] = 32'h44484000;
        data[12][34] = 32'h44488000;
        data[12][35] = 32'h4448c000;
        data[12][36] = 32'h44490000;
        data[12][37] = 32'h44494000;
        data[12][38] = 32'h44498000;
        data[12][39] = 32'h4449c000;
        data[12][40] = 32'h444a0000;
        data[12][41] = 32'h444a4000;
        data[12][42] = 32'h444a8000;
        data[12][43] = 32'h444ac000;
        data[12][44] = 32'h444b0000;
        data[12][45] = 32'h444b4000;
        data[12][46] = 32'h444b8000;
        data[12][47] = 32'h444bc000;
        data[12][48] = 32'h444c0000;
        data[12][49] = 32'h444c4000;
        data[12][50] = 32'h444c8000;
        data[12][51] = 32'h444cc000;
        data[12][52] = 32'h444d0000;
        data[12][53] = 32'h444d4000;
        data[12][54] = 32'h444d8000;
        data[12][55] = 32'h444dc000;
        data[12][56] = 32'h444e0000;
        data[12][57] = 32'h444e4000;
        data[12][58] = 32'h444e8000;
        data[12][59] = 32'h444ec000;
        data[12][60] = 32'h444f0000;
        data[12][61] = 32'h444f4000;
        data[12][62] = 32'h444f8000;
        data[12][63] = 32'h444fc000;
        data[13][0] = 32'h44500000;
        data[13][1] = 32'h44504000;
        data[13][2] = 32'h44508000;
        data[13][3] = 32'h4450c000;
        data[13][4] = 32'h44510000;
        data[13][5] = 32'h44514000;
        data[13][6] = 32'h44518000;
        data[13][7] = 32'h4451c000;
        data[13][8] = 32'h44520000;
        data[13][9] = 32'h44524000;
        data[13][10] = 32'h44528000;
        data[13][11] = 32'h4452c000;
        data[13][12] = 32'h44530000;
        data[13][13] = 32'h44534000;
        data[13][14] = 32'h44538000;
        data[13][15] = 32'h4453c000;
        data[13][16] = 32'h44540000;
        data[13][17] = 32'h44544000;
        data[13][18] = 32'h44548000;
        data[13][19] = 32'h4454c000;
        data[13][20] = 32'h44550000;
        data[13][21] = 32'h44554000;
        data[13][22] = 32'h44558000;
        data[13][23] = 32'h4455c000;
        data[13][24] = 32'h44560000;
        data[13][25] = 32'h44564000;
        data[13][26] = 32'h44568000;
        data[13][27] = 32'h4456c000;
        data[13][28] = 32'h44570000;
        data[13][29] = 32'h44574000;
        data[13][30] = 32'h44578000;
        data[13][31] = 32'h4457c000;
        data[13][32] = 32'h44580000;
        data[13][33] = 32'h44584000;
        data[13][34] = 32'h44588000;
        data[13][35] = 32'h4458c000;
        data[13][36] = 32'h44590000;
        data[13][37] = 32'h44594000;
        data[13][38] = 32'h44598000;
        data[13][39] = 32'h4459c000;
        data[13][40] = 32'h445a0000;
        data[13][41] = 32'h445a4000;
        data[13][42] = 32'h445a8000;
        data[13][43] = 32'h445ac000;
        data[13][44] = 32'h445b0000;
        data[13][45] = 32'h445b4000;
        data[13][46] = 32'h445b8000;
        data[13][47] = 32'h445bc000;
        data[13][48] = 32'h445c0000;
        data[13][49] = 32'h445c4000;
        data[13][50] = 32'h445c8000;
        data[13][51] = 32'h445cc000;
        data[13][52] = 32'h445d0000;
        data[13][53] = 32'h445d4000;
        data[13][54] = 32'h445d8000;
        data[13][55] = 32'h445dc000;
        data[13][56] = 32'h445e0000;
        data[13][57] = 32'h445e4000;
        data[13][58] = 32'h445e8000;
        data[13][59] = 32'h445ec000;
        data[13][60] = 32'h445f0000;
        data[13][61] = 32'h445f4000;
        data[13][62] = 32'h445f8000;
        data[13][63] = 32'h445fc000;
        data[14][0] = 32'h44600000;
        data[14][1] = 32'h44604000;
        data[14][2] = 32'h44608000;
        data[14][3] = 32'h4460c000;
        data[14][4] = 32'h44610000;
        data[14][5] = 32'h44614000;
        data[14][6] = 32'h44618000;
        data[14][7] = 32'h4461c000;
        data[14][8] = 32'h44620000;
        data[14][9] = 32'h44624000;
        data[14][10] = 32'h44628000;
        data[14][11] = 32'h4462c000;
        data[14][12] = 32'h44630000;
        data[14][13] = 32'h44634000;
        data[14][14] = 32'h44638000;
        data[14][15] = 32'h4463c000;
        data[14][16] = 32'h44640000;
        data[14][17] = 32'h44644000;
        data[14][18] = 32'h44648000;
        data[14][19] = 32'h4464c000;
        data[14][20] = 32'h44650000;
        data[14][21] = 32'h44654000;
        data[14][22] = 32'h44658000;
        data[14][23] = 32'h4465c000;
        data[14][24] = 32'h44660000;
        data[14][25] = 32'h44664000;
        data[14][26] = 32'h44668000;
        data[14][27] = 32'h4466c000;
        data[14][28] = 32'h44670000;
        data[14][29] = 32'h44674000;
        data[14][30] = 32'h44678000;
        data[14][31] = 32'h4467c000;
        data[14][32] = 32'h44680000;
        data[14][33] = 32'h44684000;
        data[14][34] = 32'h44688000;
        data[14][35] = 32'h4468c000;
        data[14][36] = 32'h44690000;
        data[14][37] = 32'h44694000;
        data[14][38] = 32'h44698000;
        data[14][39] = 32'h4469c000;
        data[14][40] = 32'h446a0000;
        data[14][41] = 32'h446a4000;
        data[14][42] = 32'h446a8000;
        data[14][43] = 32'h446ac000;
        data[14][44] = 32'h446b0000;
        data[14][45] = 32'h446b4000;
        data[14][46] = 32'h446b8000;
        data[14][47] = 32'h446bc000;
        data[14][48] = 32'h446c0000;
        data[14][49] = 32'h446c4000;
        data[14][50] = 32'h446c8000;
        data[14][51] = 32'h446cc000;
        data[14][52] = 32'h446d0000;
        data[14][53] = 32'h446d4000;
        data[14][54] = 32'h446d8000;
        data[14][55] = 32'h446dc000;
        data[14][56] = 32'h446e0000;
        data[14][57] = 32'h446e4000;
        data[14][58] = 32'h446e8000;
        data[14][59] = 32'h446ec000;
        data[14][60] = 32'h446f0000;
        data[14][61] = 32'h446f4000;
        data[14][62] = 32'h446f8000;
        data[14][63] = 32'h446fc000;
        data[15][0] = 32'h44700000;
        data[15][1] = 32'h44704000;
        data[15][2] = 32'h44708000;
        data[15][3] = 32'h4470c000;
        data[15][4] = 32'h44710000;
        data[15][5] = 32'h44714000;
        data[15][6] = 32'h44718000;
        data[15][7] = 32'h4471c000;
        data[15][8] = 32'h44720000;
        data[15][9] = 32'h44724000;
        data[15][10] = 32'h44728000;
        data[15][11] = 32'h4472c000;
        data[15][12] = 32'h44730000;
        data[15][13] = 32'h44734000;
        data[15][14] = 32'h44738000;
        data[15][15] = 32'h4473c000;
        data[15][16] = 32'h44740000;
        data[15][17] = 32'h44744000;
        data[15][18] = 32'h44748000;
        data[15][19] = 32'h4474c000;
        data[15][20] = 32'h44750000;
        data[15][21] = 32'h44754000;
        data[15][22] = 32'h44758000;
        data[15][23] = 32'h4475c000;
        data[15][24] = 32'h44760000;
        data[15][25] = 32'h44764000;
        data[15][26] = 32'h44768000;
        data[15][27] = 32'h4476c000;
        data[15][28] = 32'h44770000;
        data[15][29] = 32'h44774000;
        data[15][30] = 32'h44778000;
        data[15][31] = 32'h4477c000;
        data[15][32] = 32'h44780000;
        data[15][33] = 32'h44784000;
        data[15][34] = 32'h44788000;
        data[15][35] = 32'h4478c000;
        data[15][36] = 32'h44790000;
        data[15][37] = 32'h44794000;
        data[15][38] = 32'h44798000;
        data[15][39] = 32'h4479c000;
        data[15][40] = 32'h447a0000;
        data[15][41] = 32'h447a4000;
        data[15][42] = 32'h447a8000;
        data[15][43] = 32'h447ac000;
        data[15][44] = 32'h447b0000;
        data[15][45] = 32'h447b4000;
        data[15][46] = 32'h447b8000;
        data[15][47] = 32'h447bc000;
        data[15][48] = 32'h447c0000;
        data[15][49] = 32'h447c4000;
        data[15][50] = 32'h447c8000;
        data[15][51] = 32'h447cc000;
        data[15][52] = 32'h447d0000;
        data[15][53] = 32'h447d4000;
        data[15][54] = 32'h447d8000;
        data[15][55] = 32'h447dc000;
        data[15][56] = 32'h447e0000;
        data[15][57] = 32'h447e4000;
        data[15][58] = 32'h447e8000;
        data[15][59] = 32'h447ec000;
        data[15][60] = 32'h447f0000;
        data[15][61] = 32'h447f4000;
        data[15][62] = 32'h447f8000;
        data[15][63] = 32'h447fc000;
        data[16][0] = 32'h44800000;
        data[16][1] = 32'h44802000;
        data[16][2] = 32'h44804000;
        data[16][3] = 32'h44806000;
        data[16][4] = 32'h44808000;
        data[16][5] = 32'h4480a000;
        data[16][6] = 32'h4480c000;
        data[16][7] = 32'h4480e000;
        data[16][8] = 32'h44810000;
        data[16][9] = 32'h44812000;
        data[16][10] = 32'h44814000;
        data[16][11] = 32'h44816000;
        data[16][12] = 32'h44818000;
        data[16][13] = 32'h4481a000;
        data[16][14] = 32'h4481c000;
        data[16][15] = 32'h4481e000;
        data[16][16] = 32'h44820000;
        data[16][17] = 32'h44822000;
        data[16][18] = 32'h44824000;
        data[16][19] = 32'h44826000;
        data[16][20] = 32'h44828000;
        data[16][21] = 32'h4482a000;
        data[16][22] = 32'h4482c000;
        data[16][23] = 32'h4482e000;
        data[16][24] = 32'h44830000;
        data[16][25] = 32'h44832000;
        data[16][26] = 32'h44834000;
        data[16][27] = 32'h44836000;
        data[16][28] = 32'h44838000;
        data[16][29] = 32'h4483a000;
        data[16][30] = 32'h4483c000;
        data[16][31] = 32'h4483e000;
        data[16][32] = 32'h44840000;
        data[16][33] = 32'h44842000;
        data[16][34] = 32'h44844000;
        data[16][35] = 32'h44846000;
        data[16][36] = 32'h44848000;
        data[16][37] = 32'h4484a000;
        data[16][38] = 32'h4484c000;
        data[16][39] = 32'h4484e000;
        data[16][40] = 32'h44850000;
        data[16][41] = 32'h44852000;
        data[16][42] = 32'h44854000;
        data[16][43] = 32'h44856000;
        data[16][44] = 32'h44858000;
        data[16][45] = 32'h4485a000;
        data[16][46] = 32'h4485c000;
        data[16][47] = 32'h4485e000;
        data[16][48] = 32'h44860000;
        data[16][49] = 32'h44862000;
        data[16][50] = 32'h44864000;
        data[16][51] = 32'h44866000;
        data[16][52] = 32'h44868000;
        data[16][53] = 32'h4486a000;
        data[16][54] = 32'h4486c000;
        data[16][55] = 32'h4486e000;
        data[16][56] = 32'h44870000;
        data[16][57] = 32'h44872000;
        data[16][58] = 32'h44874000;
        data[16][59] = 32'h44876000;
        data[16][60] = 32'h44878000;
        data[16][61] = 32'h4487a000;
        data[16][62] = 32'h4487c000;
        data[16][63] = 32'h4487e000;
        data[17][0] = 32'h44880000;
        data[17][1] = 32'h44882000;
        data[17][2] = 32'h44884000;
        data[17][3] = 32'h44886000;
        data[17][4] = 32'h44888000;
        data[17][5] = 32'h4488a000;
        data[17][6] = 32'h4488c000;
        data[17][7] = 32'h4488e000;
        data[17][8] = 32'h44890000;
        data[17][9] = 32'h44892000;
        data[17][10] = 32'h44894000;
        data[17][11] = 32'h44896000;
        data[17][12] = 32'h44898000;
        data[17][13] = 32'h4489a000;
        data[17][14] = 32'h4489c000;
        data[17][15] = 32'h4489e000;
        data[17][16] = 32'h448a0000;
        data[17][17] = 32'h448a2000;
        data[17][18] = 32'h448a4000;
        data[17][19] = 32'h448a6000;
        data[17][20] = 32'h448a8000;
        data[17][21] = 32'h448aa000;
        data[17][22] = 32'h448ac000;
        data[17][23] = 32'h448ae000;
        data[17][24] = 32'h448b0000;
        data[17][25] = 32'h448b2000;
        data[17][26] = 32'h448b4000;
        data[17][27] = 32'h448b6000;
        data[17][28] = 32'h448b8000;
        data[17][29] = 32'h448ba000;
        data[17][30] = 32'h448bc000;
        data[17][31] = 32'h448be000;
        data[17][32] = 32'h448c0000;
        data[17][33] = 32'h448c2000;
        data[17][34] = 32'h448c4000;
        data[17][35] = 32'h448c6000;
        data[17][36] = 32'h448c8000;
        data[17][37] = 32'h448ca000;
        data[17][38] = 32'h448cc000;
        data[17][39] = 32'h448ce000;
        data[17][40] = 32'h448d0000;
        data[17][41] = 32'h448d2000;
        data[17][42] = 32'h448d4000;
        data[17][43] = 32'h448d6000;
        data[17][44] = 32'h448d8000;
        data[17][45] = 32'h448da000;
        data[17][46] = 32'h448dc000;
        data[17][47] = 32'h448de000;
        data[17][48] = 32'h448e0000;
        data[17][49] = 32'h448e2000;
        data[17][50] = 32'h448e4000;
        data[17][51] = 32'h448e6000;
        data[17][52] = 32'h448e8000;
        data[17][53] = 32'h448ea000;
        data[17][54] = 32'h448ec000;
        data[17][55] = 32'h448ee000;
        data[17][56] = 32'h448f0000;
        data[17][57] = 32'h448f2000;
        data[17][58] = 32'h448f4000;
        data[17][59] = 32'h448f6000;
        data[17][60] = 32'h448f8000;
        data[17][61] = 32'h448fa000;
        data[17][62] = 32'h448fc000;
        data[17][63] = 32'h448fe000;
        data[18][0] = 32'h44900000;
        data[18][1] = 32'h44902000;
        data[18][2] = 32'h44904000;
        data[18][3] = 32'h44906000;
        data[18][4] = 32'h44908000;
        data[18][5] = 32'h4490a000;
        data[18][6] = 32'h4490c000;
        data[18][7] = 32'h4490e000;
        data[18][8] = 32'h44910000;
        data[18][9] = 32'h44912000;
        data[18][10] = 32'h44914000;
        data[18][11] = 32'h44916000;
        data[18][12] = 32'h44918000;
        data[18][13] = 32'h4491a000;
        data[18][14] = 32'h4491c000;
        data[18][15] = 32'h4491e000;
        data[18][16] = 32'h44920000;
        data[18][17] = 32'h44922000;
        data[18][18] = 32'h44924000;
        data[18][19] = 32'h44926000;
        data[18][20] = 32'h44928000;
        data[18][21] = 32'h4492a000;
        data[18][22] = 32'h4492c000;
        data[18][23] = 32'h4492e000;
        data[18][24] = 32'h44930000;
        data[18][25] = 32'h44932000;
        data[18][26] = 32'h44934000;
        data[18][27] = 32'h44936000;
        data[18][28] = 32'h44938000;
        data[18][29] = 32'h4493a000;
        data[18][30] = 32'h4493c000;
        data[18][31] = 32'h4493e000;
        data[18][32] = 32'h44940000;
        data[18][33] = 32'h44942000;
        data[18][34] = 32'h44944000;
        data[18][35] = 32'h44946000;
        data[18][36] = 32'h44948000;
        data[18][37] = 32'h4494a000;
        data[18][38] = 32'h4494c000;
        data[18][39] = 32'h4494e000;
        data[18][40] = 32'h44950000;
        data[18][41] = 32'h44952000;
        data[18][42] = 32'h44954000;
        data[18][43] = 32'h44956000;
        data[18][44] = 32'h44958000;
        data[18][45] = 32'h4495a000;
        data[18][46] = 32'h4495c000;
        data[18][47] = 32'h4495e000;
        data[18][48] = 32'h44960000;
        data[18][49] = 32'h44962000;
        data[18][50] = 32'h44964000;
        data[18][51] = 32'h44966000;
        data[18][52] = 32'h44968000;
        data[18][53] = 32'h4496a000;
        data[18][54] = 32'h4496c000;
        data[18][55] = 32'h4496e000;
        data[18][56] = 32'h44970000;
        data[18][57] = 32'h44972000;
        data[18][58] = 32'h44974000;
        data[18][59] = 32'h44976000;
        data[18][60] = 32'h44978000;
        data[18][61] = 32'h4497a000;
        data[18][62] = 32'h4497c000;
        data[18][63] = 32'h4497e000;
        data[19][0] = 32'h44980000;
        data[19][1] = 32'h44982000;
        data[19][2] = 32'h44984000;
        data[19][3] = 32'h44986000;
        data[19][4] = 32'h44988000;
        data[19][5] = 32'h4498a000;
        data[19][6] = 32'h4498c000;
        data[19][7] = 32'h4498e000;
        data[19][8] = 32'h44990000;
        data[19][9] = 32'h44992000;
        data[19][10] = 32'h44994000;
        data[19][11] = 32'h44996000;
        data[19][12] = 32'h44998000;
        data[19][13] = 32'h4499a000;
        data[19][14] = 32'h4499c000;
        data[19][15] = 32'h4499e000;
        data[19][16] = 32'h449a0000;
        data[19][17] = 32'h449a2000;
        data[19][18] = 32'h449a4000;
        data[19][19] = 32'h449a6000;
        data[19][20] = 32'h449a8000;
        data[19][21] = 32'h449aa000;
        data[19][22] = 32'h449ac000;
        data[19][23] = 32'h449ae000;
        data[19][24] = 32'h449b0000;
        data[19][25] = 32'h449b2000;
        data[19][26] = 32'h449b4000;
        data[19][27] = 32'h449b6000;
        data[19][28] = 32'h449b8000;
        data[19][29] = 32'h449ba000;
        data[19][30] = 32'h449bc000;
        data[19][31] = 32'h449be000;
        data[19][32] = 32'h449c0000;
        data[19][33] = 32'h449c2000;
        data[19][34] = 32'h449c4000;
        data[19][35] = 32'h449c6000;
        data[19][36] = 32'h449c8000;
        data[19][37] = 32'h449ca000;
        data[19][38] = 32'h449cc000;
        data[19][39] = 32'h449ce000;
        data[19][40] = 32'h449d0000;
        data[19][41] = 32'h449d2000;
        data[19][42] = 32'h449d4000;
        data[19][43] = 32'h449d6000;
        data[19][44] = 32'h449d8000;
        data[19][45] = 32'h449da000;
        data[19][46] = 32'h449dc000;
        data[19][47] = 32'h449de000;
        data[19][48] = 32'h449e0000;
        data[19][49] = 32'h449e2000;
        data[19][50] = 32'h449e4000;
        data[19][51] = 32'h449e6000;
        data[19][52] = 32'h449e8000;
        data[19][53] = 32'h449ea000;
        data[19][54] = 32'h449ec000;
        data[19][55] = 32'h449ee000;
        data[19][56] = 32'h449f0000;
        data[19][57] = 32'h449f2000;
        data[19][58] = 32'h449f4000;
        data[19][59] = 32'h449f6000;
        data[19][60] = 32'h449f8000;
        data[19][61] = 32'h449fa000;
        data[19][62] = 32'h449fc000;
        data[19][63] = 32'h449fe000;
        data[20][0] = 32'h44a00000;
        data[20][1] = 32'h44a02000;
        data[20][2] = 32'h44a04000;
        data[20][3] = 32'h44a06000;
        data[20][4] = 32'h44a08000;
        data[20][5] = 32'h44a0a000;
        data[20][6] = 32'h44a0c000;
        data[20][7] = 32'h44a0e000;
        data[20][8] = 32'h44a10000;
        data[20][9] = 32'h44a12000;
        data[20][10] = 32'h44a14000;
        data[20][11] = 32'h44a16000;
        data[20][12] = 32'h44a18000;
        data[20][13] = 32'h44a1a000;
        data[20][14] = 32'h44a1c000;
        data[20][15] = 32'h44a1e000;
        data[20][16] = 32'h44a20000;
        data[20][17] = 32'h44a22000;
        data[20][18] = 32'h44a24000;
        data[20][19] = 32'h44a26000;
        data[20][20] = 32'h44a28000;
        data[20][21] = 32'h44a2a000;
        data[20][22] = 32'h44a2c000;
        data[20][23] = 32'h44a2e000;
        data[20][24] = 32'h44a30000;
        data[20][25] = 32'h44a32000;
        data[20][26] = 32'h44a34000;
        data[20][27] = 32'h44a36000;
        data[20][28] = 32'h44a38000;
        data[20][29] = 32'h44a3a000;
        data[20][30] = 32'h44a3c000;
        data[20][31] = 32'h44a3e000;
        data[20][32] = 32'h44a40000;
        data[20][33] = 32'h44a42000;
        data[20][34] = 32'h44a44000;
        data[20][35] = 32'h44a46000;
        data[20][36] = 32'h44a48000;
        data[20][37] = 32'h44a4a000;
        data[20][38] = 32'h44a4c000;
        data[20][39] = 32'h44a4e000;
        data[20][40] = 32'h44a50000;
        data[20][41] = 32'h44a52000;
        data[20][42] = 32'h44a54000;
        data[20][43] = 32'h44a56000;
        data[20][44] = 32'h44a58000;
        data[20][45] = 32'h44a5a000;
        data[20][46] = 32'h44a5c000;
        data[20][47] = 32'h44a5e000;
        data[20][48] = 32'h44a60000;
        data[20][49] = 32'h44a62000;
        data[20][50] = 32'h44a64000;
        data[20][51] = 32'h44a66000;
        data[20][52] = 32'h44a68000;
        data[20][53] = 32'h44a6a000;
        data[20][54] = 32'h44a6c000;
        data[20][55] = 32'h44a6e000;
        data[20][56] = 32'h44a70000;
        data[20][57] = 32'h44a72000;
        data[20][58] = 32'h44a74000;
        data[20][59] = 32'h44a76000;
        data[20][60] = 32'h44a78000;
        data[20][61] = 32'h44a7a000;
        data[20][62] = 32'h44a7c000;
        data[20][63] = 32'h44a7e000;
        data[21][0] = 32'h44a80000;
        data[21][1] = 32'h44a82000;
        data[21][2] = 32'h44a84000;
        data[21][3] = 32'h44a86000;
        data[21][4] = 32'h44a88000;
        data[21][5] = 32'h44a8a000;
        data[21][6] = 32'h44a8c000;
        data[21][7] = 32'h44a8e000;
        data[21][8] = 32'h44a90000;
        data[21][9] = 32'h44a92000;
        data[21][10] = 32'h44a94000;
        data[21][11] = 32'h44a96000;
        data[21][12] = 32'h44a98000;
        data[21][13] = 32'h44a9a000;
        data[21][14] = 32'h44a9c000;
        data[21][15] = 32'h44a9e000;
        data[21][16] = 32'h44aa0000;
        data[21][17] = 32'h44aa2000;
        data[21][18] = 32'h44aa4000;
        data[21][19] = 32'h44aa6000;
        data[21][20] = 32'h44aa8000;
        data[21][21] = 32'h44aaa000;
        data[21][22] = 32'h44aac000;
        data[21][23] = 32'h44aae000;
        data[21][24] = 32'h44ab0000;
        data[21][25] = 32'h44ab2000;
        data[21][26] = 32'h44ab4000;
        data[21][27] = 32'h44ab6000;
        data[21][28] = 32'h44ab8000;
        data[21][29] = 32'h44aba000;
        data[21][30] = 32'h44abc000;
        data[21][31] = 32'h44abe000;
        data[21][32] = 32'h44ac0000;
        data[21][33] = 32'h44ac2000;
        data[21][34] = 32'h44ac4000;
        data[21][35] = 32'h44ac6000;
        data[21][36] = 32'h44ac8000;
        data[21][37] = 32'h44aca000;
        data[21][38] = 32'h44acc000;
        data[21][39] = 32'h44ace000;
        data[21][40] = 32'h44ad0000;
        data[21][41] = 32'h44ad2000;
        data[21][42] = 32'h44ad4000;
        data[21][43] = 32'h44ad6000;
        data[21][44] = 32'h44ad8000;
        data[21][45] = 32'h44ada000;
        data[21][46] = 32'h44adc000;
        data[21][47] = 32'h44ade000;
        data[21][48] = 32'h44ae0000;
        data[21][49] = 32'h44ae2000;
        data[21][50] = 32'h44ae4000;
        data[21][51] = 32'h44ae6000;
        data[21][52] = 32'h44ae8000;
        data[21][53] = 32'h44aea000;
        data[21][54] = 32'h44aec000;
        data[21][55] = 32'h44aee000;
        data[21][56] = 32'h44af0000;
        data[21][57] = 32'h44af2000;
        data[21][58] = 32'h44af4000;
        data[21][59] = 32'h44af6000;
        data[21][60] = 32'h44af8000;
        data[21][61] = 32'h44afa000;
        data[21][62] = 32'h44afc000;
        data[21][63] = 32'h44afe000;
        data[22][0] = 32'h44b00000;
        data[22][1] = 32'h44b02000;
        data[22][2] = 32'h44b04000;
        data[22][3] = 32'h44b06000;
        data[22][4] = 32'h44b08000;
        data[22][5] = 32'h44b0a000;
        data[22][6] = 32'h44b0c000;
        data[22][7] = 32'h44b0e000;
        data[22][8] = 32'h44b10000;
        data[22][9] = 32'h44b12000;
        data[22][10] = 32'h44b14000;
        data[22][11] = 32'h44b16000;
        data[22][12] = 32'h44b18000;
        data[22][13] = 32'h44b1a000;
        data[22][14] = 32'h44b1c000;
        data[22][15] = 32'h44b1e000;
        data[22][16] = 32'h44b20000;
        data[22][17] = 32'h44b22000;
        data[22][18] = 32'h44b24000;
        data[22][19] = 32'h44b26000;
        data[22][20] = 32'h44b28000;
        data[22][21] = 32'h44b2a000;
        data[22][22] = 32'h44b2c000;
        data[22][23] = 32'h44b2e000;
        data[22][24] = 32'h44b30000;
        data[22][25] = 32'h44b32000;
        data[22][26] = 32'h44b34000;
        data[22][27] = 32'h44b36000;
        data[22][28] = 32'h44b38000;
        data[22][29] = 32'h44b3a000;
        data[22][30] = 32'h44b3c000;
        data[22][31] = 32'h44b3e000;
        data[22][32] = 32'h44b40000;
        data[22][33] = 32'h44b42000;
        data[22][34] = 32'h44b44000;
        data[22][35] = 32'h44b46000;
        data[22][36] = 32'h44b48000;
        data[22][37] = 32'h44b4a000;
        data[22][38] = 32'h44b4c000;
        data[22][39] = 32'h44b4e000;
        data[22][40] = 32'h44b50000;
        data[22][41] = 32'h44b52000;
        data[22][42] = 32'h44b54000;
        data[22][43] = 32'h44b56000;
        data[22][44] = 32'h44b58000;
        data[22][45] = 32'h44b5a000;
        data[22][46] = 32'h44b5c000;
        data[22][47] = 32'h44b5e000;
        data[22][48] = 32'h44b60000;
        data[22][49] = 32'h44b62000;
        data[22][50] = 32'h44b64000;
        data[22][51] = 32'h44b66000;
        data[22][52] = 32'h44b68000;
        data[22][53] = 32'h44b6a000;
        data[22][54] = 32'h44b6c000;
        data[22][55] = 32'h44b6e000;
        data[22][56] = 32'h44b70000;
        data[22][57] = 32'h44b72000;
        data[22][58] = 32'h44b74000;
        data[22][59] = 32'h44b76000;
        data[22][60] = 32'h44b78000;
        data[22][61] = 32'h44b7a000;
        data[22][62] = 32'h44b7c000;
        data[22][63] = 32'h44b7e000;
        data[23][0] = 32'h44b80000;
        data[23][1] = 32'h44b82000;
        data[23][2] = 32'h44b84000;
        data[23][3] = 32'h44b86000;
        data[23][4] = 32'h44b88000;
        data[23][5] = 32'h44b8a000;
        data[23][6] = 32'h44b8c000;
        data[23][7] = 32'h44b8e000;
        data[23][8] = 32'h44b90000;
        data[23][9] = 32'h44b92000;
        data[23][10] = 32'h44b94000;
        data[23][11] = 32'h44b96000;
        data[23][12] = 32'h44b98000;
        data[23][13] = 32'h44b9a000;
        data[23][14] = 32'h44b9c000;
        data[23][15] = 32'h44b9e000;
        data[23][16] = 32'h44ba0000;
        data[23][17] = 32'h44ba2000;
        data[23][18] = 32'h44ba4000;
        data[23][19] = 32'h44ba6000;
        data[23][20] = 32'h44ba8000;
        data[23][21] = 32'h44baa000;
        data[23][22] = 32'h44bac000;
        data[23][23] = 32'h44bae000;
        data[23][24] = 32'h44bb0000;
        data[23][25] = 32'h44bb2000;
        data[23][26] = 32'h44bb4000;
        data[23][27] = 32'h44bb6000;
        data[23][28] = 32'h44bb8000;
        data[23][29] = 32'h44bba000;
        data[23][30] = 32'h44bbc000;
        data[23][31] = 32'h44bbe000;
        data[23][32] = 32'h44bc0000;
        data[23][33] = 32'h44bc2000;
        data[23][34] = 32'h44bc4000;
        data[23][35] = 32'h44bc6000;
        data[23][36] = 32'h44bc8000;
        data[23][37] = 32'h44bca000;
        data[23][38] = 32'h44bcc000;
        data[23][39] = 32'h44bce000;
        data[23][40] = 32'h44bd0000;
        data[23][41] = 32'h44bd2000;
        data[23][42] = 32'h44bd4000;
        data[23][43] = 32'h44bd6000;
        data[23][44] = 32'h44bd8000;
        data[23][45] = 32'h44bda000;
        data[23][46] = 32'h44bdc000;
        data[23][47] = 32'h44bde000;
        data[23][48] = 32'h44be0000;
        data[23][49] = 32'h44be2000;
        data[23][50] = 32'h44be4000;
        data[23][51] = 32'h44be6000;
        data[23][52] = 32'h44be8000;
        data[23][53] = 32'h44bea000;
        data[23][54] = 32'h44bec000;
        data[23][55] = 32'h44bee000;
        data[23][56] = 32'h44bf0000;
        data[23][57] = 32'h44bf2000;
        data[23][58] = 32'h44bf4000;
        data[23][59] = 32'h44bf6000;
        data[23][60] = 32'h44bf8000;
        data[23][61] = 32'h44bfa000;
        data[23][62] = 32'h44bfc000;
        data[23][63] = 32'h44bfe000;
        data[24][0] = 32'h44c00000;
        data[24][1] = 32'h44c02000;
        data[24][2] = 32'h44c04000;
        data[24][3] = 32'h44c06000;
        data[24][4] = 32'h44c08000;
        data[24][5] = 32'h44c0a000;
        data[24][6] = 32'h44c0c000;
        data[24][7] = 32'h44c0e000;
        data[24][8] = 32'h44c10000;
        data[24][9] = 32'h44c12000;
        data[24][10] = 32'h44c14000;
        data[24][11] = 32'h44c16000;
        data[24][12] = 32'h44c18000;
        data[24][13] = 32'h44c1a000;
        data[24][14] = 32'h44c1c000;
        data[24][15] = 32'h44c1e000;
        data[24][16] = 32'h44c20000;
        data[24][17] = 32'h44c22000;
        data[24][18] = 32'h44c24000;
        data[24][19] = 32'h44c26000;
        data[24][20] = 32'h44c28000;
        data[24][21] = 32'h44c2a000;
        data[24][22] = 32'h44c2c000;
        data[24][23] = 32'h44c2e000;
        data[24][24] = 32'h44c30000;
        data[24][25] = 32'h44c32000;
        data[24][26] = 32'h44c34000;
        data[24][27] = 32'h44c36000;
        data[24][28] = 32'h44c38000;
        data[24][29] = 32'h44c3a000;
        data[24][30] = 32'h44c3c000;
        data[24][31] = 32'h44c3e000;
        data[24][32] = 32'h44c40000;
        data[24][33] = 32'h44c42000;
        data[24][34] = 32'h44c44000;
        data[24][35] = 32'h44c46000;
        data[24][36] = 32'h44c48000;
        data[24][37] = 32'h44c4a000;
        data[24][38] = 32'h44c4c000;
        data[24][39] = 32'h44c4e000;
        data[24][40] = 32'h44c50000;
        data[24][41] = 32'h44c52000;
        data[24][42] = 32'h44c54000;
        data[24][43] = 32'h44c56000;
        data[24][44] = 32'h44c58000;
        data[24][45] = 32'h44c5a000;
        data[24][46] = 32'h44c5c000;
        data[24][47] = 32'h44c5e000;
        data[24][48] = 32'h44c60000;
        data[24][49] = 32'h44c62000;
        data[24][50] = 32'h44c64000;
        data[24][51] = 32'h44c66000;
        data[24][52] = 32'h44c68000;
        data[24][53] = 32'h44c6a000;
        data[24][54] = 32'h44c6c000;
        data[24][55] = 32'h44c6e000;
        data[24][56] = 32'h44c70000;
        data[24][57] = 32'h44c72000;
        data[24][58] = 32'h44c74000;
        data[24][59] = 32'h44c76000;
        data[24][60] = 32'h44c78000;
        data[24][61] = 32'h44c7a000;
        data[24][62] = 32'h44c7c000;
        data[24][63] = 32'h44c7e000;
        data[25][0] = 32'h44c80000;
        data[25][1] = 32'h44c82000;
        data[25][2] = 32'h44c84000;
        data[25][3] = 32'h44c86000;
        data[25][4] = 32'h44c88000;
        data[25][5] = 32'h44c8a000;
        data[25][6] = 32'h44c8c000;
        data[25][7] = 32'h44c8e000;
        data[25][8] = 32'h44c90000;
        data[25][9] = 32'h44c92000;
        data[25][10] = 32'h44c94000;
        data[25][11] = 32'h44c96000;
        data[25][12] = 32'h44c98000;
        data[25][13] = 32'h44c9a000;
        data[25][14] = 32'h44c9c000;
        data[25][15] = 32'h44c9e000;
        data[25][16] = 32'h44ca0000;
        data[25][17] = 32'h44ca2000;
        data[25][18] = 32'h44ca4000;
        data[25][19] = 32'h44ca6000;
        data[25][20] = 32'h44ca8000;
        data[25][21] = 32'h44caa000;
        data[25][22] = 32'h44cac000;
        data[25][23] = 32'h44cae000;
        data[25][24] = 32'h44cb0000;
        data[25][25] = 32'h44cb2000;
        data[25][26] = 32'h44cb4000;
        data[25][27] = 32'h44cb6000;
        data[25][28] = 32'h44cb8000;
        data[25][29] = 32'h44cba000;
        data[25][30] = 32'h44cbc000;
        data[25][31] = 32'h44cbe000;
        data[25][32] = 32'h44cc0000;
        data[25][33] = 32'h44cc2000;
        data[25][34] = 32'h44cc4000;
        data[25][35] = 32'h44cc6000;
        data[25][36] = 32'h44cc8000;
        data[25][37] = 32'h44cca000;
        data[25][38] = 32'h44ccc000;
        data[25][39] = 32'h44cce000;
        data[25][40] = 32'h44cd0000;
        data[25][41] = 32'h44cd2000;
        data[25][42] = 32'h44cd4000;
        data[25][43] = 32'h44cd6000;
        data[25][44] = 32'h44cd8000;
        data[25][45] = 32'h44cda000;
        data[25][46] = 32'h44cdc000;
        data[25][47] = 32'h44cde000;
        data[25][48] = 32'h44ce0000;
        data[25][49] = 32'h44ce2000;
        data[25][50] = 32'h44ce4000;
        data[25][51] = 32'h44ce6000;
        data[25][52] = 32'h44ce8000;
        data[25][53] = 32'h44cea000;
        data[25][54] = 32'h44cec000;
        data[25][55] = 32'h44cee000;
        data[25][56] = 32'h44cf0000;
        data[25][57] = 32'h44cf2000;
        data[25][58] = 32'h44cf4000;
        data[25][59] = 32'h44cf6000;
        data[25][60] = 32'h44cf8000;
        data[25][61] = 32'h44cfa000;
        data[25][62] = 32'h44cfc000;
        data[25][63] = 32'h44cfe000;
        data[26][0] = 32'h44d00000;
        data[26][1] = 32'h44d02000;
        data[26][2] = 32'h44d04000;
        data[26][3] = 32'h44d06000;
        data[26][4] = 32'h44d08000;
        data[26][5] = 32'h44d0a000;
        data[26][6] = 32'h44d0c000;
        data[26][7] = 32'h44d0e000;
        data[26][8] = 32'h44d10000;
        data[26][9] = 32'h44d12000;
        data[26][10] = 32'h44d14000;
        data[26][11] = 32'h44d16000;
        data[26][12] = 32'h44d18000;
        data[26][13] = 32'h44d1a000;
        data[26][14] = 32'h44d1c000;
        data[26][15] = 32'h44d1e000;
        data[26][16] = 32'h44d20000;
        data[26][17] = 32'h44d22000;
        data[26][18] = 32'h44d24000;
        data[26][19] = 32'h44d26000;
        data[26][20] = 32'h44d28000;
        data[26][21] = 32'h44d2a000;
        data[26][22] = 32'h44d2c000;
        data[26][23] = 32'h44d2e000;
        data[26][24] = 32'h44d30000;
        data[26][25] = 32'h44d32000;
        data[26][26] = 32'h44d34000;
        data[26][27] = 32'h44d36000;
        data[26][28] = 32'h44d38000;
        data[26][29] = 32'h44d3a000;
        data[26][30] = 32'h44d3c000;
        data[26][31] = 32'h44d3e000;
        data[26][32] = 32'h44d40000;
        data[26][33] = 32'h44d42000;
        data[26][34] = 32'h44d44000;
        data[26][35] = 32'h44d46000;
        data[26][36] = 32'h44d48000;
        data[26][37] = 32'h44d4a000;
        data[26][38] = 32'h44d4c000;
        data[26][39] = 32'h44d4e000;
        data[26][40] = 32'h44d50000;
        data[26][41] = 32'h44d52000;
        data[26][42] = 32'h44d54000;
        data[26][43] = 32'h44d56000;
        data[26][44] = 32'h44d58000;
        data[26][45] = 32'h44d5a000;
        data[26][46] = 32'h44d5c000;
        data[26][47] = 32'h44d5e000;
        data[26][48] = 32'h44d60000;
        data[26][49] = 32'h44d62000;
        data[26][50] = 32'h44d64000;
        data[26][51] = 32'h44d66000;
        data[26][52] = 32'h44d68000;
        data[26][53] = 32'h44d6a000;
        data[26][54] = 32'h44d6c000;
        data[26][55] = 32'h44d6e000;
        data[26][56] = 32'h44d70000;
        data[26][57] = 32'h44d72000;
        data[26][58] = 32'h44d74000;
        data[26][59] = 32'h44d76000;
        data[26][60] = 32'h44d78000;
        data[26][61] = 32'h44d7a000;
        data[26][62] = 32'h44d7c000;
        data[26][63] = 32'h44d7e000;
        data[27][0] = 32'h44d80000;
        data[27][1] = 32'h44d82000;
        data[27][2] = 32'h44d84000;
        data[27][3] = 32'h44d86000;
        data[27][4] = 32'h44d88000;
        data[27][5] = 32'h44d8a000;
        data[27][6] = 32'h44d8c000;
        data[27][7] = 32'h44d8e000;
        data[27][8] = 32'h44d90000;
        data[27][9] = 32'h44d92000;
        data[27][10] = 32'h44d94000;
        data[27][11] = 32'h44d96000;
        data[27][12] = 32'h44d98000;
        data[27][13] = 32'h44d9a000;
        data[27][14] = 32'h44d9c000;
        data[27][15] = 32'h44d9e000;
        data[27][16] = 32'h44da0000;
        data[27][17] = 32'h44da2000;
        data[27][18] = 32'h44da4000;
        data[27][19] = 32'h44da6000;
        data[27][20] = 32'h44da8000;
        data[27][21] = 32'h44daa000;
        data[27][22] = 32'h44dac000;
        data[27][23] = 32'h44dae000;
        data[27][24] = 32'h44db0000;
        data[27][25] = 32'h44db2000;
        data[27][26] = 32'h44db4000;
        data[27][27] = 32'h44db6000;
        data[27][28] = 32'h44db8000;
        data[27][29] = 32'h44dba000;
        data[27][30] = 32'h44dbc000;
        data[27][31] = 32'h44dbe000;
        data[27][32] = 32'h44dc0000;
        data[27][33] = 32'h44dc2000;
        data[27][34] = 32'h44dc4000;
        data[27][35] = 32'h44dc6000;
        data[27][36] = 32'h44dc8000;
        data[27][37] = 32'h44dca000;
        data[27][38] = 32'h44dcc000;
        data[27][39] = 32'h44dce000;
        data[27][40] = 32'h44dd0000;
        data[27][41] = 32'h44dd2000;
        data[27][42] = 32'h44dd4000;
        data[27][43] = 32'h44dd6000;
        data[27][44] = 32'h44dd8000;
        data[27][45] = 32'h44dda000;
        data[27][46] = 32'h44ddc000;
        data[27][47] = 32'h44dde000;
        data[27][48] = 32'h44de0000;
        data[27][49] = 32'h44de2000;
        data[27][50] = 32'h44de4000;
        data[27][51] = 32'h44de6000;
        data[27][52] = 32'h44de8000;
        data[27][53] = 32'h44dea000;
        data[27][54] = 32'h44dec000;
        data[27][55] = 32'h44dee000;
        data[27][56] = 32'h44df0000;
        data[27][57] = 32'h44df2000;
        data[27][58] = 32'h44df4000;
        data[27][59] = 32'h44df6000;
        data[27][60] = 32'h44df8000;
        data[27][61] = 32'h44dfa000;
        data[27][62] = 32'h44dfc000;
        data[27][63] = 32'h44dfe000;
        data[28][0] = 32'h44e00000;
        data[28][1] = 32'h44e02000;
        data[28][2] = 32'h44e04000;
        data[28][3] = 32'h44e06000;
        data[28][4] = 32'h44e08000;
        data[28][5] = 32'h44e0a000;
        data[28][6] = 32'h44e0c000;
        data[28][7] = 32'h44e0e000;
        data[28][8] = 32'h44e10000;
        data[28][9] = 32'h44e12000;
        data[28][10] = 32'h44e14000;
        data[28][11] = 32'h44e16000;
        data[28][12] = 32'h44e18000;
        data[28][13] = 32'h44e1a000;
        data[28][14] = 32'h44e1c000;
        data[28][15] = 32'h44e1e000;
        data[28][16] = 32'h44e20000;
        data[28][17] = 32'h44e22000;
        data[28][18] = 32'h44e24000;
        data[28][19] = 32'h44e26000;
        data[28][20] = 32'h44e28000;
        data[28][21] = 32'h44e2a000;
        data[28][22] = 32'h44e2c000;
        data[28][23] = 32'h44e2e000;
        data[28][24] = 32'h44e30000;
        data[28][25] = 32'h44e32000;
        data[28][26] = 32'h44e34000;
        data[28][27] = 32'h44e36000;
        data[28][28] = 32'h44e38000;
        data[28][29] = 32'h44e3a000;
        data[28][30] = 32'h44e3c000;
        data[28][31] = 32'h44e3e000;
        data[28][32] = 32'h44e40000;
        data[28][33] = 32'h44e42000;
        data[28][34] = 32'h44e44000;
        data[28][35] = 32'h44e46000;
        data[28][36] = 32'h44e48000;
        data[28][37] = 32'h44e4a000;
        data[28][38] = 32'h44e4c000;
        data[28][39] = 32'h44e4e000;
        data[28][40] = 32'h44e50000;
        data[28][41] = 32'h44e52000;
        data[28][42] = 32'h44e54000;
        data[28][43] = 32'h44e56000;
        data[28][44] = 32'h44e58000;
        data[28][45] = 32'h44e5a000;
        data[28][46] = 32'h44e5c000;
        data[28][47] = 32'h44e5e000;
        data[28][48] = 32'h44e60000;
        data[28][49] = 32'h44e62000;
        data[28][50] = 32'h44e64000;
        data[28][51] = 32'h44e66000;
        data[28][52] = 32'h44e68000;
        data[28][53] = 32'h44e6a000;
        data[28][54] = 32'h44e6c000;
        data[28][55] = 32'h44e6e000;
        data[28][56] = 32'h44e70000;
        data[28][57] = 32'h44e72000;
        data[28][58] = 32'h44e74000;
        data[28][59] = 32'h44e76000;
        data[28][60] = 32'h44e78000;
        data[28][61] = 32'h44e7a000;
        data[28][62] = 32'h44e7c000;
        data[28][63] = 32'h44e7e000;
        data[29][0] = 32'h44e80000;
        data[29][1] = 32'h44e82000;
        data[29][2] = 32'h44e84000;
        data[29][3] = 32'h44e86000;
        data[29][4] = 32'h44e88000;
        data[29][5] = 32'h44e8a000;
        data[29][6] = 32'h44e8c000;
        data[29][7] = 32'h44e8e000;
        data[29][8] = 32'h44e90000;
        data[29][9] = 32'h44e92000;
        data[29][10] = 32'h44e94000;
        data[29][11] = 32'h44e96000;
        data[29][12] = 32'h44e98000;
        data[29][13] = 32'h44e9a000;
        data[29][14] = 32'h44e9c000;
        data[29][15] = 32'h44e9e000;
        data[29][16] = 32'h44ea0000;
        data[29][17] = 32'h44ea2000;
        data[29][18] = 32'h44ea4000;
        data[29][19] = 32'h44ea6000;
        data[29][20] = 32'h44ea8000;
        data[29][21] = 32'h44eaa000;
        data[29][22] = 32'h44eac000;
        data[29][23] = 32'h44eae000;
        data[29][24] = 32'h44eb0000;
        data[29][25] = 32'h44eb2000;
        data[29][26] = 32'h44eb4000;
        data[29][27] = 32'h44eb6000;
        data[29][28] = 32'h44eb8000;
        data[29][29] = 32'h44eba000;
        data[29][30] = 32'h44ebc000;
        data[29][31] = 32'h44ebe000;
        data[29][32] = 32'h44ec0000;
        data[29][33] = 32'h44ec2000;
        data[29][34] = 32'h44ec4000;
        data[29][35] = 32'h44ec6000;
        data[29][36] = 32'h44ec8000;
        data[29][37] = 32'h44eca000;
        data[29][38] = 32'h44ecc000;
        data[29][39] = 32'h44ece000;
        data[29][40] = 32'h44ed0000;
        data[29][41] = 32'h44ed2000;
        data[29][42] = 32'h44ed4000;
        data[29][43] = 32'h44ed6000;
        data[29][44] = 32'h44ed8000;
        data[29][45] = 32'h44eda000;
        data[29][46] = 32'h44edc000;
        data[29][47] = 32'h44ede000;
        data[29][48] = 32'h44ee0000;
        data[29][49] = 32'h44ee2000;
        data[29][50] = 32'h44ee4000;
        data[29][51] = 32'h44ee6000;
        data[29][52] = 32'h44ee8000;
        data[29][53] = 32'h44eea000;
        data[29][54] = 32'h44eec000;
        data[29][55] = 32'h44eee000;
        data[29][56] = 32'h44ef0000;
        data[29][57] = 32'h44ef2000;
        data[29][58] = 32'h44ef4000;
        data[29][59] = 32'h44ef6000;
        data[29][60] = 32'h44ef8000;
        data[29][61] = 32'h44efa000;
        data[29][62] = 32'h44efc000;
        data[29][63] = 32'h44efe000;
        data[30][0] = 32'h44f00000;
        data[30][1] = 32'h44f02000;
        data[30][2] = 32'h44f04000;
        data[30][3] = 32'h44f06000;
        data[30][4] = 32'h44f08000;
        data[30][5] = 32'h44f0a000;
        data[30][6] = 32'h44f0c000;
        data[30][7] = 32'h44f0e000;
        data[30][8] = 32'h44f10000;
        data[30][9] = 32'h44f12000;
        data[30][10] = 32'h44f14000;
        data[30][11] = 32'h44f16000;
        data[30][12] = 32'h44f18000;
        data[30][13] = 32'h44f1a000;
        data[30][14] = 32'h44f1c000;
        data[30][15] = 32'h44f1e000;
        data[30][16] = 32'h44f20000;
        data[30][17] = 32'h44f22000;
        data[30][18] = 32'h44f24000;
        data[30][19] = 32'h44f26000;
        data[30][20] = 32'h44f28000;
        data[30][21] = 32'h44f2a000;
        data[30][22] = 32'h44f2c000;
        data[30][23] = 32'h44f2e000;
        data[30][24] = 32'h44f30000;
        data[30][25] = 32'h44f32000;
        data[30][26] = 32'h44f34000;
        data[30][27] = 32'h44f36000;
        data[30][28] = 32'h44f38000;
        data[30][29] = 32'h44f3a000;
        data[30][30] = 32'h44f3c000;
        data[30][31] = 32'h44f3e000;
        data[30][32] = 32'h44f40000;
        data[30][33] = 32'h44f42000;
        data[30][34] = 32'h44f44000;
        data[30][35] = 32'h44f46000;
        data[30][36] = 32'h44f48000;
        data[30][37] = 32'h44f4a000;
        data[30][38] = 32'h44f4c000;
        data[30][39] = 32'h44f4e000;
        data[30][40] = 32'h44f50000;
        data[30][41] = 32'h44f52000;
        data[30][42] = 32'h44f54000;
        data[30][43] = 32'h44f56000;
        data[30][44] = 32'h44f58000;
        data[30][45] = 32'h44f5a000;
        data[30][46] = 32'h44f5c000;
        data[30][47] = 32'h44f5e000;
        data[30][48] = 32'h44f60000;
        data[30][49] = 32'h44f62000;
        data[30][50] = 32'h44f64000;
        data[30][51] = 32'h44f66000;
        data[30][52] = 32'h44f68000;
        data[30][53] = 32'h44f6a000;
        data[30][54] = 32'h44f6c000;
        data[30][55] = 32'h44f6e000;
        data[30][56] = 32'h44f70000;
        data[30][57] = 32'h44f72000;
        data[30][58] = 32'h44f74000;
        data[30][59] = 32'h44f76000;
        data[30][60] = 32'h44f78000;
        data[30][61] = 32'h44f7a000;
        data[30][62] = 32'h44f7c000;
        data[30][63] = 32'h44f7e000;
        data[31][0] = 32'h44f80000;
        data[31][1] = 32'h44f82000;
        data[31][2] = 32'h44f84000;
        data[31][3] = 32'h44f86000;
        data[31][4] = 32'h44f88000;
        data[31][5] = 32'h44f8a000;
        data[31][6] = 32'h44f8c000;
        data[31][7] = 32'h44f8e000;
        data[31][8] = 32'h44f90000;
        data[31][9] = 32'h44f92000;
        data[31][10] = 32'h44f94000;
        data[31][11] = 32'h44f96000;
        data[31][12] = 32'h44f98000;
        data[31][13] = 32'h44f9a000;
        data[31][14] = 32'h44f9c000;
        data[31][15] = 32'h44f9e000;
        data[31][16] = 32'h44fa0000;
        data[31][17] = 32'h44fa2000;
        data[31][18] = 32'h44fa4000;
        data[31][19] = 32'h44fa6000;
        data[31][20] = 32'h44fa8000;
        data[31][21] = 32'h44faa000;
        data[31][22] = 32'h44fac000;
        data[31][23] = 32'h44fae000;
        data[31][24] = 32'h44fb0000;
        data[31][25] = 32'h44fb2000;
        data[31][26] = 32'h44fb4000;
        data[31][27] = 32'h44fb6000;
        data[31][28] = 32'h44fb8000;
        data[31][29] = 32'h44fba000;
        data[31][30] = 32'h44fbc000;
        data[31][31] = 32'h44fbe000;
        data[31][32] = 32'h44fc0000;
        data[31][33] = 32'h44fc2000;
        data[31][34] = 32'h44fc4000;
        data[31][35] = 32'h44fc6000;
        data[31][36] = 32'h44fc8000;
        data[31][37] = 32'h44fca000;
        data[31][38] = 32'h44fcc000;
        data[31][39] = 32'h44fce000;
        data[31][40] = 32'h44fd0000;
        data[31][41] = 32'h44fd2000;
        data[31][42] = 32'h44fd4000;
        data[31][43] = 32'h44fd6000;
        data[31][44] = 32'h44fd8000;
        data[31][45] = 32'h44fda000;
        data[31][46] = 32'h44fdc000;
        data[31][47] = 32'h44fde000;
        data[31][48] = 32'h44fe0000;
        data[31][49] = 32'h44fe2000;
        data[31][50] = 32'h44fe4000;
        data[31][51] = 32'h44fe6000;
        data[31][52] = 32'h44fe8000;
        data[31][53] = 32'h44fea000;
        data[31][54] = 32'h44fec000;
        data[31][55] = 32'h44fee000;
        data[31][56] = 32'h44ff0000;
        data[31][57] = 32'h44ff2000;
        data[31][58] = 32'h44ff4000;
        data[31][59] = 32'h44ff6000;
        data[31][60] = 32'h44ff8000;
        data[31][61] = 32'h44ffa000;
        data[31][62] = 32'h44ffc000;
        data[31][63] = 32'h44ffe000;
        data[32][0] = 32'h45000000;
        data[32][1] = 32'h45001000;
        data[32][2] = 32'h45002000;
        data[32][3] = 32'h45003000;
        data[32][4] = 32'h45004000;
        data[32][5] = 32'h45005000;
        data[32][6] = 32'h45006000;
        data[32][7] = 32'h45007000;
        data[32][8] = 32'h45008000;
        data[32][9] = 32'h45009000;
        data[32][10] = 32'h4500a000;
        data[32][11] = 32'h4500b000;
        data[32][12] = 32'h4500c000;
        data[32][13] = 32'h4500d000;
        data[32][14] = 32'h4500e000;
        data[32][15] = 32'h4500f000;
        data[32][16] = 32'h45010000;
        data[32][17] = 32'h45011000;
        data[32][18] = 32'h45012000;
        data[32][19] = 32'h45013000;
        data[32][20] = 32'h45014000;
        data[32][21] = 32'h45015000;
        data[32][22] = 32'h45016000;
        data[32][23] = 32'h45017000;
        data[32][24] = 32'h45018000;
        data[32][25] = 32'h45019000;
        data[32][26] = 32'h4501a000;
        data[32][27] = 32'h4501b000;
        data[32][28] = 32'h4501c000;
        data[32][29] = 32'h4501d000;
        data[32][30] = 32'h4501e000;
        data[32][31] = 32'h4501f000;
        data[32][32] = 32'h45020000;
        data[32][33] = 32'h45021000;
        data[32][34] = 32'h45022000;
        data[32][35] = 32'h45023000;
        data[32][36] = 32'h45024000;
        data[32][37] = 32'h45025000;
        data[32][38] = 32'h45026000;
        data[32][39] = 32'h45027000;
        data[32][40] = 32'h45028000;
        data[32][41] = 32'h45029000;
        data[32][42] = 32'h4502a000;
        data[32][43] = 32'h4502b000;
        data[32][44] = 32'h4502c000;
        data[32][45] = 32'h4502d000;
        data[32][46] = 32'h4502e000;
        data[32][47] = 32'h4502f000;
        data[32][48] = 32'h45030000;
        data[32][49] = 32'h45031000;
        data[32][50] = 32'h45032000;
        data[32][51] = 32'h45033000;
        data[32][52] = 32'h45034000;
        data[32][53] = 32'h45035000;
        data[32][54] = 32'h45036000;
        data[32][55] = 32'h45037000;
        data[32][56] = 32'h45038000;
        data[32][57] = 32'h45039000;
        data[32][58] = 32'h4503a000;
        data[32][59] = 32'h4503b000;
        data[32][60] = 32'h4503c000;
        data[32][61] = 32'h4503d000;
        data[32][62] = 32'h4503e000;
        data[32][63] = 32'h4503f000;
        data[33][0] = 32'h45040000;
        data[33][1] = 32'h45041000;
        data[33][2] = 32'h45042000;
        data[33][3] = 32'h45043000;
        data[33][4] = 32'h45044000;
        data[33][5] = 32'h45045000;
        data[33][6] = 32'h45046000;
        data[33][7] = 32'h45047000;
        data[33][8] = 32'h45048000;
        data[33][9] = 32'h45049000;
        data[33][10] = 32'h4504a000;
        data[33][11] = 32'h4504b000;
        data[33][12] = 32'h4504c000;
        data[33][13] = 32'h4504d000;
        data[33][14] = 32'h4504e000;
        data[33][15] = 32'h4504f000;
        data[33][16] = 32'h45050000;
        data[33][17] = 32'h45051000;
        data[33][18] = 32'h45052000;
        data[33][19] = 32'h45053000;
        data[33][20] = 32'h45054000;
        data[33][21] = 32'h45055000;
        data[33][22] = 32'h45056000;
        data[33][23] = 32'h45057000;
        data[33][24] = 32'h45058000;
        data[33][25] = 32'h45059000;
        data[33][26] = 32'h4505a000;
        data[33][27] = 32'h4505b000;
        data[33][28] = 32'h4505c000;
        data[33][29] = 32'h4505d000;
        data[33][30] = 32'h4505e000;
        data[33][31] = 32'h4505f000;
        data[33][32] = 32'h45060000;
        data[33][33] = 32'h45061000;
        data[33][34] = 32'h45062000;
        data[33][35] = 32'h45063000;
        data[33][36] = 32'h45064000;
        data[33][37] = 32'h45065000;
        data[33][38] = 32'h45066000;
        data[33][39] = 32'h45067000;
        data[33][40] = 32'h45068000;
        data[33][41] = 32'h45069000;
        data[33][42] = 32'h4506a000;
        data[33][43] = 32'h4506b000;
        data[33][44] = 32'h4506c000;
        data[33][45] = 32'h4506d000;
        data[33][46] = 32'h4506e000;
        data[33][47] = 32'h4506f000;
        data[33][48] = 32'h45070000;
        data[33][49] = 32'h45071000;
        data[33][50] = 32'h45072000;
        data[33][51] = 32'h45073000;
        data[33][52] = 32'h45074000;
        data[33][53] = 32'h45075000;
        data[33][54] = 32'h45076000;
        data[33][55] = 32'h45077000;
        data[33][56] = 32'h45078000;
        data[33][57] = 32'h45079000;
        data[33][58] = 32'h4507a000;
        data[33][59] = 32'h4507b000;
        data[33][60] = 32'h4507c000;
        data[33][61] = 32'h4507d000;
        data[33][62] = 32'h4507e000;
        data[33][63] = 32'h4507f000;
        data[34][0] = 32'h45080000;
        data[34][1] = 32'h45081000;
        data[34][2] = 32'h45082000;
        data[34][3] = 32'h45083000;
        data[34][4] = 32'h45084000;
        data[34][5] = 32'h45085000;
        data[34][6] = 32'h45086000;
        data[34][7] = 32'h45087000;
        data[34][8] = 32'h45088000;
        data[34][9] = 32'h45089000;
        data[34][10] = 32'h4508a000;
        data[34][11] = 32'h4508b000;
        data[34][12] = 32'h4508c000;
        data[34][13] = 32'h4508d000;
        data[34][14] = 32'h4508e000;
        data[34][15] = 32'h4508f000;
        data[34][16] = 32'h45090000;
        data[34][17] = 32'h45091000;
        data[34][18] = 32'h45092000;
        data[34][19] = 32'h45093000;
        data[34][20] = 32'h45094000;
        data[34][21] = 32'h45095000;
        data[34][22] = 32'h45096000;
        data[34][23] = 32'h45097000;
        data[34][24] = 32'h45098000;
        data[34][25] = 32'h45099000;
        data[34][26] = 32'h4509a000;
        data[34][27] = 32'h4509b000;
        data[34][28] = 32'h4509c000;
        data[34][29] = 32'h4509d000;
        data[34][30] = 32'h4509e000;
        data[34][31] = 32'h4509f000;
        data[34][32] = 32'h450a0000;
        data[34][33] = 32'h450a1000;
        data[34][34] = 32'h450a2000;
        data[34][35] = 32'h450a3000;
        data[34][36] = 32'h450a4000;
        data[34][37] = 32'h450a5000;
        data[34][38] = 32'h450a6000;
        data[34][39] = 32'h450a7000;
        data[34][40] = 32'h450a8000;
        data[34][41] = 32'h450a9000;
        data[34][42] = 32'h450aa000;
        data[34][43] = 32'h450ab000;
        data[34][44] = 32'h450ac000;
        data[34][45] = 32'h450ad000;
        data[34][46] = 32'h450ae000;
        data[34][47] = 32'h450af000;
        data[34][48] = 32'h450b0000;
        data[34][49] = 32'h450b1000;
        data[34][50] = 32'h450b2000;
        data[34][51] = 32'h450b3000;
        data[34][52] = 32'h450b4000;
        data[34][53] = 32'h450b5000;
        data[34][54] = 32'h450b6000;
        data[34][55] = 32'h450b7000;
        data[34][56] = 32'h450b8000;
        data[34][57] = 32'h450b9000;
        data[34][58] = 32'h450ba000;
        data[34][59] = 32'h450bb000;
        data[34][60] = 32'h450bc000;
        data[34][61] = 32'h450bd000;
        data[34][62] = 32'h450be000;
        data[34][63] = 32'h450bf000;
        data[35][0] = 32'h450c0000;
        data[35][1] = 32'h450c1000;
        data[35][2] = 32'h450c2000;
        data[35][3] = 32'h450c3000;
        data[35][4] = 32'h450c4000;
        data[35][5] = 32'h450c5000;
        data[35][6] = 32'h450c6000;
        data[35][7] = 32'h450c7000;
        data[35][8] = 32'h450c8000;
        data[35][9] = 32'h450c9000;
        data[35][10] = 32'h450ca000;
        data[35][11] = 32'h450cb000;
        data[35][12] = 32'h450cc000;
        data[35][13] = 32'h450cd000;
        data[35][14] = 32'h450ce000;
        data[35][15] = 32'h450cf000;
        data[35][16] = 32'h450d0000;
        data[35][17] = 32'h450d1000;
        data[35][18] = 32'h450d2000;
        data[35][19] = 32'h450d3000;
        data[35][20] = 32'h450d4000;
        data[35][21] = 32'h450d5000;
        data[35][22] = 32'h450d6000;
        data[35][23] = 32'h450d7000;
        data[35][24] = 32'h450d8000;
        data[35][25] = 32'h450d9000;
        data[35][26] = 32'h450da000;
        data[35][27] = 32'h450db000;
        data[35][28] = 32'h450dc000;
        data[35][29] = 32'h450dd000;
        data[35][30] = 32'h450de000;
        data[35][31] = 32'h450df000;
        data[35][32] = 32'h450e0000;
        data[35][33] = 32'h450e1000;
        data[35][34] = 32'h450e2000;
        data[35][35] = 32'h450e3000;
        data[35][36] = 32'h450e4000;
        data[35][37] = 32'h450e5000;
        data[35][38] = 32'h450e6000;
        data[35][39] = 32'h450e7000;
        data[35][40] = 32'h450e8000;
        data[35][41] = 32'h450e9000;
        data[35][42] = 32'h450ea000;
        data[35][43] = 32'h450eb000;
        data[35][44] = 32'h450ec000;
        data[35][45] = 32'h450ed000;
        data[35][46] = 32'h450ee000;
        data[35][47] = 32'h450ef000;
        data[35][48] = 32'h450f0000;
        data[35][49] = 32'h450f1000;
        data[35][50] = 32'h450f2000;
        data[35][51] = 32'h450f3000;
        data[35][52] = 32'h450f4000;
        data[35][53] = 32'h450f5000;
        data[35][54] = 32'h450f6000;
        data[35][55] = 32'h450f7000;
        data[35][56] = 32'h450f8000;
        data[35][57] = 32'h450f9000;
        data[35][58] = 32'h450fa000;
        data[35][59] = 32'h450fb000;
        data[35][60] = 32'h450fc000;
        data[35][61] = 32'h450fd000;
        data[35][62] = 32'h450fe000;
        data[35][63] = 32'h450ff000;
        data[36][0] = 32'h45100000;
        data[36][1] = 32'h45101000;
        data[36][2] = 32'h45102000;
        data[36][3] = 32'h45103000;
        data[36][4] = 32'h45104000;
        data[36][5] = 32'h45105000;
        data[36][6] = 32'h45106000;
        data[36][7] = 32'h45107000;
        data[36][8] = 32'h45108000;
        data[36][9] = 32'h45109000;
        data[36][10] = 32'h4510a000;
        data[36][11] = 32'h4510b000;
        data[36][12] = 32'h4510c000;
        data[36][13] = 32'h4510d000;
        data[36][14] = 32'h4510e000;
        data[36][15] = 32'h4510f000;
        data[36][16] = 32'h45110000;
        data[36][17] = 32'h45111000;
        data[36][18] = 32'h45112000;
        data[36][19] = 32'h45113000;
        data[36][20] = 32'h45114000;
        data[36][21] = 32'h45115000;
        data[36][22] = 32'h45116000;
        data[36][23] = 32'h45117000;
        data[36][24] = 32'h45118000;
        data[36][25] = 32'h45119000;
        data[36][26] = 32'h4511a000;
        data[36][27] = 32'h4511b000;
        data[36][28] = 32'h4511c000;
        data[36][29] = 32'h4511d000;
        data[36][30] = 32'h4511e000;
        data[36][31] = 32'h4511f000;
        data[36][32] = 32'h45120000;
        data[36][33] = 32'h45121000;
        data[36][34] = 32'h45122000;
        data[36][35] = 32'h45123000;
        data[36][36] = 32'h45124000;
        data[36][37] = 32'h45125000;
        data[36][38] = 32'h45126000;
        data[36][39] = 32'h45127000;
        data[36][40] = 32'h45128000;
        data[36][41] = 32'h45129000;
        data[36][42] = 32'h4512a000;
        data[36][43] = 32'h4512b000;
        data[36][44] = 32'h4512c000;
        data[36][45] = 32'h4512d000;
        data[36][46] = 32'h4512e000;
        data[36][47] = 32'h4512f000;
        data[36][48] = 32'h45130000;
        data[36][49] = 32'h45131000;
        data[36][50] = 32'h45132000;
        data[36][51] = 32'h45133000;
        data[36][52] = 32'h45134000;
        data[36][53] = 32'h45135000;
        data[36][54] = 32'h45136000;
        data[36][55] = 32'h45137000;
        data[36][56] = 32'h45138000;
        data[36][57] = 32'h45139000;
        data[36][58] = 32'h4513a000;
        data[36][59] = 32'h4513b000;
        data[36][60] = 32'h4513c000;
        data[36][61] = 32'h4513d000;
        data[36][62] = 32'h4513e000;
        data[36][63] = 32'h4513f000;
        data[37][0] = 32'h45140000;
        data[37][1] = 32'h45141000;
        data[37][2] = 32'h45142000;
        data[37][3] = 32'h45143000;
        data[37][4] = 32'h45144000;
        data[37][5] = 32'h45145000;
        data[37][6] = 32'h45146000;
        data[37][7] = 32'h45147000;
        data[37][8] = 32'h45148000;
        data[37][9] = 32'h45149000;
        data[37][10] = 32'h4514a000;
        data[37][11] = 32'h4514b000;
        data[37][12] = 32'h4514c000;
        data[37][13] = 32'h4514d000;
        data[37][14] = 32'h4514e000;
        data[37][15] = 32'h4514f000;
        data[37][16] = 32'h45150000;
        data[37][17] = 32'h45151000;
        data[37][18] = 32'h45152000;
        data[37][19] = 32'h45153000;
        data[37][20] = 32'h45154000;
        data[37][21] = 32'h45155000;
        data[37][22] = 32'h45156000;
        data[37][23] = 32'h45157000;
        data[37][24] = 32'h45158000;
        data[37][25] = 32'h45159000;
        data[37][26] = 32'h4515a000;
        data[37][27] = 32'h4515b000;
        data[37][28] = 32'h4515c000;
        data[37][29] = 32'h4515d000;
        data[37][30] = 32'h4515e000;
        data[37][31] = 32'h4515f000;
        data[37][32] = 32'h45160000;
        data[37][33] = 32'h45161000;
        data[37][34] = 32'h45162000;
        data[37][35] = 32'h45163000;
        data[37][36] = 32'h45164000;
        data[37][37] = 32'h45165000;
        data[37][38] = 32'h45166000;
        data[37][39] = 32'h45167000;
        data[37][40] = 32'h45168000;
        data[37][41] = 32'h45169000;
        data[37][42] = 32'h4516a000;
        data[37][43] = 32'h4516b000;
        data[37][44] = 32'h4516c000;
        data[37][45] = 32'h4516d000;
        data[37][46] = 32'h4516e000;
        data[37][47] = 32'h4516f000;
        data[37][48] = 32'h45170000;
        data[37][49] = 32'h45171000;
        data[37][50] = 32'h45172000;
        data[37][51] = 32'h45173000;
        data[37][52] = 32'h45174000;
        data[37][53] = 32'h45175000;
        data[37][54] = 32'h45176000;
        data[37][55] = 32'h45177000;
        data[37][56] = 32'h45178000;
        data[37][57] = 32'h45179000;
        data[37][58] = 32'h4517a000;
        data[37][59] = 32'h4517b000;
        data[37][60] = 32'h4517c000;
        data[37][61] = 32'h4517d000;
        data[37][62] = 32'h4517e000;
        data[37][63] = 32'h4517f000;
        data[38][0] = 32'h45180000;
        data[38][1] = 32'h45181000;
        data[38][2] = 32'h45182000;
        data[38][3] = 32'h45183000;
        data[38][4] = 32'h45184000;
        data[38][5] = 32'h45185000;
        data[38][6] = 32'h45186000;
        data[38][7] = 32'h45187000;
        data[38][8] = 32'h45188000;
        data[38][9] = 32'h45189000;
        data[38][10] = 32'h4518a000;
        data[38][11] = 32'h4518b000;
        data[38][12] = 32'h4518c000;
        data[38][13] = 32'h4518d000;
        data[38][14] = 32'h4518e000;
        data[38][15] = 32'h4518f000;
        data[38][16] = 32'h45190000;
        data[38][17] = 32'h45191000;
        data[38][18] = 32'h45192000;
        data[38][19] = 32'h45193000;
        data[38][20] = 32'h45194000;
        data[38][21] = 32'h45195000;
        data[38][22] = 32'h45196000;
        data[38][23] = 32'h45197000;
        data[38][24] = 32'h45198000;
        data[38][25] = 32'h45199000;
        data[38][26] = 32'h4519a000;
        data[38][27] = 32'h4519b000;
        data[38][28] = 32'h4519c000;
        data[38][29] = 32'h4519d000;
        data[38][30] = 32'h4519e000;
        data[38][31] = 32'h4519f000;
        data[38][32] = 32'h451a0000;
        data[38][33] = 32'h451a1000;
        data[38][34] = 32'h451a2000;
        data[38][35] = 32'h451a3000;
        data[38][36] = 32'h451a4000;
        data[38][37] = 32'h451a5000;
        data[38][38] = 32'h451a6000;
        data[38][39] = 32'h451a7000;
        data[38][40] = 32'h451a8000;
        data[38][41] = 32'h451a9000;
        data[38][42] = 32'h451aa000;
        data[38][43] = 32'h451ab000;
        data[38][44] = 32'h451ac000;
        data[38][45] = 32'h451ad000;
        data[38][46] = 32'h451ae000;
        data[38][47] = 32'h451af000;
        data[38][48] = 32'h451b0000;
        data[38][49] = 32'h451b1000;
        data[38][50] = 32'h451b2000;
        data[38][51] = 32'h451b3000;
        data[38][52] = 32'h451b4000;
        data[38][53] = 32'h451b5000;
        data[38][54] = 32'h451b6000;
        data[38][55] = 32'h451b7000;
        data[38][56] = 32'h451b8000;
        data[38][57] = 32'h451b9000;
        data[38][58] = 32'h451ba000;
        data[38][59] = 32'h451bb000;
        data[38][60] = 32'h451bc000;
        data[38][61] = 32'h451bd000;
        data[38][62] = 32'h451be000;
        data[38][63] = 32'h451bf000;
        data[39][0] = 32'h451c0000;
        data[39][1] = 32'h451c1000;
        data[39][2] = 32'h451c2000;
        data[39][3] = 32'h451c3000;
        data[39][4] = 32'h451c4000;
        data[39][5] = 32'h451c5000;
        data[39][6] = 32'h451c6000;
        data[39][7] = 32'h451c7000;
        data[39][8] = 32'h451c8000;
        data[39][9] = 32'h451c9000;
        data[39][10] = 32'h451ca000;
        data[39][11] = 32'h451cb000;
        data[39][12] = 32'h451cc000;
        data[39][13] = 32'h451cd000;
        data[39][14] = 32'h451ce000;
        data[39][15] = 32'h451cf000;
        data[39][16] = 32'h451d0000;
        data[39][17] = 32'h451d1000;
        data[39][18] = 32'h451d2000;
        data[39][19] = 32'h451d3000;
        data[39][20] = 32'h451d4000;
        data[39][21] = 32'h451d5000;
        data[39][22] = 32'h451d6000;
        data[39][23] = 32'h451d7000;
        data[39][24] = 32'h451d8000;
        data[39][25] = 32'h451d9000;
        data[39][26] = 32'h451da000;
        data[39][27] = 32'h451db000;
        data[39][28] = 32'h451dc000;
        data[39][29] = 32'h451dd000;
        data[39][30] = 32'h451de000;
        data[39][31] = 32'h451df000;
        data[39][32] = 32'h451e0000;
        data[39][33] = 32'h451e1000;
        data[39][34] = 32'h451e2000;
        data[39][35] = 32'h451e3000;
        data[39][36] = 32'h451e4000;
        data[39][37] = 32'h451e5000;
        data[39][38] = 32'h451e6000;
        data[39][39] = 32'h451e7000;
        data[39][40] = 32'h451e8000;
        data[39][41] = 32'h451e9000;
        data[39][42] = 32'h451ea000;
        data[39][43] = 32'h451eb000;
        data[39][44] = 32'h451ec000;
        data[39][45] = 32'h451ed000;
        data[39][46] = 32'h451ee000;
        data[39][47] = 32'h451ef000;
        data[39][48] = 32'h451f0000;
        data[39][49] = 32'h451f1000;
        data[39][50] = 32'h451f2000;
        data[39][51] = 32'h451f3000;
        data[39][52] = 32'h451f4000;
        data[39][53] = 32'h451f5000;
        data[39][54] = 32'h451f6000;
        data[39][55] = 32'h451f7000;
        data[39][56] = 32'h451f8000;
        data[39][57] = 32'h451f9000;
        data[39][58] = 32'h451fa000;
        data[39][59] = 32'h451fb000;
        data[39][60] = 32'h451fc000;
        data[39][61] = 32'h451fd000;
        data[39][62] = 32'h451fe000;
        data[39][63] = 32'h451ff000;
        data[40][0] = 32'h45200000;
        data[40][1] = 32'h45201000;
        data[40][2] = 32'h45202000;
        data[40][3] = 32'h45203000;
        data[40][4] = 32'h45204000;
        data[40][5] = 32'h45205000;
        data[40][6] = 32'h45206000;
        data[40][7] = 32'h45207000;
        data[40][8] = 32'h45208000;
        data[40][9] = 32'h45209000;
        data[40][10] = 32'h4520a000;
        data[40][11] = 32'h4520b000;
        data[40][12] = 32'h4520c000;
        data[40][13] = 32'h4520d000;
        data[40][14] = 32'h4520e000;
        data[40][15] = 32'h4520f000;
        data[40][16] = 32'h45210000;
        data[40][17] = 32'h45211000;
        data[40][18] = 32'h45212000;
        data[40][19] = 32'h45213000;
        data[40][20] = 32'h45214000;
        data[40][21] = 32'h45215000;
        data[40][22] = 32'h45216000;
        data[40][23] = 32'h45217000;
        data[40][24] = 32'h45218000;
        data[40][25] = 32'h45219000;
        data[40][26] = 32'h4521a000;
        data[40][27] = 32'h4521b000;
        data[40][28] = 32'h4521c000;
        data[40][29] = 32'h4521d000;
        data[40][30] = 32'h4521e000;
        data[40][31] = 32'h4521f000;
        data[40][32] = 32'h45220000;
        data[40][33] = 32'h45221000;
        data[40][34] = 32'h45222000;
        data[40][35] = 32'h45223000;
        data[40][36] = 32'h45224000;
        data[40][37] = 32'h45225000;
        data[40][38] = 32'h45226000;
        data[40][39] = 32'h45227000;
        data[40][40] = 32'h45228000;
        data[40][41] = 32'h45229000;
        data[40][42] = 32'h4522a000;
        data[40][43] = 32'h4522b000;
        data[40][44] = 32'h4522c000;
        data[40][45] = 32'h4522d000;
        data[40][46] = 32'h4522e000;
        data[40][47] = 32'h4522f000;
        data[40][48] = 32'h45230000;
        data[40][49] = 32'h45231000;
        data[40][50] = 32'h45232000;
        data[40][51] = 32'h45233000;
        data[40][52] = 32'h45234000;
        data[40][53] = 32'h45235000;
        data[40][54] = 32'h45236000;
        data[40][55] = 32'h45237000;
        data[40][56] = 32'h45238000;
        data[40][57] = 32'h45239000;
        data[40][58] = 32'h4523a000;
        data[40][59] = 32'h4523b000;
        data[40][60] = 32'h4523c000;
        data[40][61] = 32'h4523d000;
        data[40][62] = 32'h4523e000;
        data[40][63] = 32'h4523f000;
        data[41][0] = 32'h45240000;
        data[41][1] = 32'h45241000;
        data[41][2] = 32'h45242000;
        data[41][3] = 32'h45243000;
        data[41][4] = 32'h45244000;
        data[41][5] = 32'h45245000;
        data[41][6] = 32'h45246000;
        data[41][7] = 32'h45247000;
        data[41][8] = 32'h45248000;
        data[41][9] = 32'h45249000;
        data[41][10] = 32'h4524a000;
        data[41][11] = 32'h4524b000;
        data[41][12] = 32'h4524c000;
        data[41][13] = 32'h4524d000;
        data[41][14] = 32'h4524e000;
        data[41][15] = 32'h4524f000;
        data[41][16] = 32'h45250000;
        data[41][17] = 32'h45251000;
        data[41][18] = 32'h45252000;
        data[41][19] = 32'h45253000;
        data[41][20] = 32'h45254000;
        data[41][21] = 32'h45255000;
        data[41][22] = 32'h45256000;
        data[41][23] = 32'h45257000;
        data[41][24] = 32'h45258000;
        data[41][25] = 32'h45259000;
        data[41][26] = 32'h4525a000;
        data[41][27] = 32'h4525b000;
        data[41][28] = 32'h4525c000;
        data[41][29] = 32'h4525d000;
        data[41][30] = 32'h4525e000;
        data[41][31] = 32'h4525f000;
        data[41][32] = 32'h45260000;
        data[41][33] = 32'h45261000;
        data[41][34] = 32'h45262000;
        data[41][35] = 32'h45263000;
        data[41][36] = 32'h45264000;
        data[41][37] = 32'h45265000;
        data[41][38] = 32'h45266000;
        data[41][39] = 32'h45267000;
        data[41][40] = 32'h45268000;
        data[41][41] = 32'h45269000;
        data[41][42] = 32'h4526a000;
        data[41][43] = 32'h4526b000;
        data[41][44] = 32'h4526c000;
        data[41][45] = 32'h4526d000;
        data[41][46] = 32'h4526e000;
        data[41][47] = 32'h4526f000;
        data[41][48] = 32'h45270000;
        data[41][49] = 32'h45271000;
        data[41][50] = 32'h45272000;
        data[41][51] = 32'h45273000;
        data[41][52] = 32'h45274000;
        data[41][53] = 32'h45275000;
        data[41][54] = 32'h45276000;
        data[41][55] = 32'h45277000;
        data[41][56] = 32'h45278000;
        data[41][57] = 32'h45279000;
        data[41][58] = 32'h4527a000;
        data[41][59] = 32'h4527b000;
        data[41][60] = 32'h4527c000;
        data[41][61] = 32'h4527d000;
        data[41][62] = 32'h4527e000;
        data[41][63] = 32'h4527f000;
        data[42][0] = 32'h45280000;
        data[42][1] = 32'h45281000;
        data[42][2] = 32'h45282000;
        data[42][3] = 32'h45283000;
        data[42][4] = 32'h45284000;
        data[42][5] = 32'h45285000;
        data[42][6] = 32'h45286000;
        data[42][7] = 32'h45287000;
        data[42][8] = 32'h45288000;
        data[42][9] = 32'h45289000;
        data[42][10] = 32'h4528a000;
        data[42][11] = 32'h4528b000;
        data[42][12] = 32'h4528c000;
        data[42][13] = 32'h4528d000;
        data[42][14] = 32'h4528e000;
        data[42][15] = 32'h4528f000;
        data[42][16] = 32'h45290000;
        data[42][17] = 32'h45291000;
        data[42][18] = 32'h45292000;
        data[42][19] = 32'h45293000;
        data[42][20] = 32'h45294000;
        data[42][21] = 32'h45295000;
        data[42][22] = 32'h45296000;
        data[42][23] = 32'h45297000;
        data[42][24] = 32'h45298000;
        data[42][25] = 32'h45299000;
        data[42][26] = 32'h4529a000;
        data[42][27] = 32'h4529b000;
        data[42][28] = 32'h4529c000;
        data[42][29] = 32'h4529d000;
        data[42][30] = 32'h4529e000;
        data[42][31] = 32'h4529f000;
        data[42][32] = 32'h452a0000;
        data[42][33] = 32'h452a1000;
        data[42][34] = 32'h452a2000;
        data[42][35] = 32'h452a3000;
        data[42][36] = 32'h452a4000;
        data[42][37] = 32'h452a5000;
        data[42][38] = 32'h452a6000;
        data[42][39] = 32'h452a7000;
        data[42][40] = 32'h452a8000;
        data[42][41] = 32'h452a9000;
        data[42][42] = 32'h452aa000;
        data[42][43] = 32'h452ab000;
        data[42][44] = 32'h452ac000;
        data[42][45] = 32'h452ad000;
        data[42][46] = 32'h452ae000;
        data[42][47] = 32'h452af000;
        data[42][48] = 32'h452b0000;
        data[42][49] = 32'h452b1000;
        data[42][50] = 32'h452b2000;
        data[42][51] = 32'h452b3000;
        data[42][52] = 32'h452b4000;
        data[42][53] = 32'h452b5000;
        data[42][54] = 32'h452b6000;
        data[42][55] = 32'h452b7000;
        data[42][56] = 32'h452b8000;
        data[42][57] = 32'h452b9000;
        data[42][58] = 32'h452ba000;
        data[42][59] = 32'h452bb000;
        data[42][60] = 32'h452bc000;
        data[42][61] = 32'h452bd000;
        data[42][62] = 32'h452be000;
        data[42][63] = 32'h452bf000;
        data[43][0] = 32'h452c0000;
        data[43][1] = 32'h452c1000;
        data[43][2] = 32'h452c2000;
        data[43][3] = 32'h452c3000;
        data[43][4] = 32'h452c4000;
        data[43][5] = 32'h452c5000;
        data[43][6] = 32'h452c6000;
        data[43][7] = 32'h452c7000;
        data[43][8] = 32'h452c8000;
        data[43][9] = 32'h452c9000;
        data[43][10] = 32'h452ca000;
        data[43][11] = 32'h452cb000;
        data[43][12] = 32'h452cc000;
        data[43][13] = 32'h452cd000;
        data[43][14] = 32'h452ce000;
        data[43][15] = 32'h452cf000;
        data[43][16] = 32'h452d0000;
        data[43][17] = 32'h452d1000;
        data[43][18] = 32'h452d2000;
        data[43][19] = 32'h452d3000;
        data[43][20] = 32'h452d4000;
        data[43][21] = 32'h452d5000;
        data[43][22] = 32'h452d6000;
        data[43][23] = 32'h452d7000;
        data[43][24] = 32'h452d8000;
        data[43][25] = 32'h452d9000;
        data[43][26] = 32'h452da000;
        data[43][27] = 32'h452db000;
        data[43][28] = 32'h452dc000;
        data[43][29] = 32'h452dd000;
        data[43][30] = 32'h452de000;
        data[43][31] = 32'h452df000;
        data[43][32] = 32'h452e0000;
        data[43][33] = 32'h452e1000;
        data[43][34] = 32'h452e2000;
        data[43][35] = 32'h452e3000;
        data[43][36] = 32'h452e4000;
        data[43][37] = 32'h452e5000;
        data[43][38] = 32'h452e6000;
        data[43][39] = 32'h452e7000;
        data[43][40] = 32'h452e8000;
        data[43][41] = 32'h452e9000;
        data[43][42] = 32'h452ea000;
        data[43][43] = 32'h452eb000;
        data[43][44] = 32'h452ec000;
        data[43][45] = 32'h452ed000;
        data[43][46] = 32'h452ee000;
        data[43][47] = 32'h452ef000;
        data[43][48] = 32'h452f0000;
        data[43][49] = 32'h452f1000;
        data[43][50] = 32'h452f2000;
        data[43][51] = 32'h452f3000;
        data[43][52] = 32'h452f4000;
        data[43][53] = 32'h452f5000;
        data[43][54] = 32'h452f6000;
        data[43][55] = 32'h452f7000;
        data[43][56] = 32'h452f8000;
        data[43][57] = 32'h452f9000;
        data[43][58] = 32'h452fa000;
        data[43][59] = 32'h452fb000;
        data[43][60] = 32'h452fc000;
        data[43][61] = 32'h452fd000;
        data[43][62] = 32'h452fe000;
        data[43][63] = 32'h452ff000;
        data[44][0] = 32'h45300000;
        data[44][1] = 32'h45301000;
        data[44][2] = 32'h45302000;
        data[44][3] = 32'h45303000;
        data[44][4] = 32'h45304000;
        data[44][5] = 32'h45305000;
        data[44][6] = 32'h45306000;
        data[44][7] = 32'h45307000;
        data[44][8] = 32'h45308000;
        data[44][9] = 32'h45309000;
        data[44][10] = 32'h4530a000;
        data[44][11] = 32'h4530b000;
        data[44][12] = 32'h4530c000;
        data[44][13] = 32'h4530d000;
        data[44][14] = 32'h4530e000;
        data[44][15] = 32'h4530f000;
        data[44][16] = 32'h45310000;
        data[44][17] = 32'h45311000;
        data[44][18] = 32'h45312000;
        data[44][19] = 32'h45313000;
        data[44][20] = 32'h45314000;
        data[44][21] = 32'h45315000;
        data[44][22] = 32'h45316000;
        data[44][23] = 32'h45317000;
        data[44][24] = 32'h45318000;
        data[44][25] = 32'h45319000;
        data[44][26] = 32'h4531a000;
        data[44][27] = 32'h4531b000;
        data[44][28] = 32'h4531c000;
        data[44][29] = 32'h4531d000;
        data[44][30] = 32'h4531e000;
        data[44][31] = 32'h4531f000;
        data[44][32] = 32'h45320000;
        data[44][33] = 32'h45321000;
        data[44][34] = 32'h45322000;
        data[44][35] = 32'h45323000;
        data[44][36] = 32'h45324000;
        data[44][37] = 32'h45325000;
        data[44][38] = 32'h45326000;
        data[44][39] = 32'h45327000;
        data[44][40] = 32'h45328000;
        data[44][41] = 32'h45329000;
        data[44][42] = 32'h4532a000;
        data[44][43] = 32'h4532b000;
        data[44][44] = 32'h4532c000;
        data[44][45] = 32'h4532d000;
        data[44][46] = 32'h4532e000;
        data[44][47] = 32'h4532f000;
        data[44][48] = 32'h45330000;
        data[44][49] = 32'h45331000;
        data[44][50] = 32'h45332000;
        data[44][51] = 32'h45333000;
        data[44][52] = 32'h45334000;
        data[44][53] = 32'h45335000;
        data[44][54] = 32'h45336000;
        data[44][55] = 32'h45337000;
        data[44][56] = 32'h45338000;
        data[44][57] = 32'h45339000;
        data[44][58] = 32'h4533a000;
        data[44][59] = 32'h4533b000;
        data[44][60] = 32'h4533c000;
        data[44][61] = 32'h4533d000;
        data[44][62] = 32'h4533e000;
        data[44][63] = 32'h4533f000;
        data[45][0] = 32'h45340000;
        data[45][1] = 32'h45341000;
        data[45][2] = 32'h45342000;
        data[45][3] = 32'h45343000;
        data[45][4] = 32'h45344000;
        data[45][5] = 32'h45345000;
        data[45][6] = 32'h45346000;
        data[45][7] = 32'h45347000;
        data[45][8] = 32'h45348000;
        data[45][9] = 32'h45349000;
        data[45][10] = 32'h4534a000;
        data[45][11] = 32'h4534b000;
        data[45][12] = 32'h4534c000;
        data[45][13] = 32'h4534d000;
        data[45][14] = 32'h4534e000;
        data[45][15] = 32'h4534f000;
        data[45][16] = 32'h45350000;
        data[45][17] = 32'h45351000;
        data[45][18] = 32'h45352000;
        data[45][19] = 32'h45353000;
        data[45][20] = 32'h45354000;
        data[45][21] = 32'h45355000;
        data[45][22] = 32'h45356000;
        data[45][23] = 32'h45357000;
        data[45][24] = 32'h45358000;
        data[45][25] = 32'h45359000;
        data[45][26] = 32'h4535a000;
        data[45][27] = 32'h4535b000;
        data[45][28] = 32'h4535c000;
        data[45][29] = 32'h4535d000;
        data[45][30] = 32'h4535e000;
        data[45][31] = 32'h4535f000;
        data[45][32] = 32'h45360000;
        data[45][33] = 32'h45361000;
        data[45][34] = 32'h45362000;
        data[45][35] = 32'h45363000;
        data[45][36] = 32'h45364000;
        data[45][37] = 32'h45365000;
        data[45][38] = 32'h45366000;
        data[45][39] = 32'h45367000;
        data[45][40] = 32'h45368000;
        data[45][41] = 32'h45369000;
        data[45][42] = 32'h4536a000;
        data[45][43] = 32'h4536b000;
        data[45][44] = 32'h4536c000;
        data[45][45] = 32'h4536d000;
        data[45][46] = 32'h4536e000;
        data[45][47] = 32'h4536f000;
        data[45][48] = 32'h45370000;
        data[45][49] = 32'h45371000;
        data[45][50] = 32'h45372000;
        data[45][51] = 32'h45373000;
        data[45][52] = 32'h45374000;
        data[45][53] = 32'h45375000;
        data[45][54] = 32'h45376000;
        data[45][55] = 32'h45377000;
        data[45][56] = 32'h45378000;
        data[45][57] = 32'h45379000;
        data[45][58] = 32'h4537a000;
        data[45][59] = 32'h4537b000;
        data[45][60] = 32'h4537c000;
        data[45][61] = 32'h4537d000;
        data[45][62] = 32'h4537e000;
        data[45][63] = 32'h4537f000;
        data[46][0] = 32'h45380000;
        data[46][1] = 32'h45381000;
        data[46][2] = 32'h45382000;
        data[46][3] = 32'h45383000;
        data[46][4] = 32'h45384000;
        data[46][5] = 32'h45385000;
        data[46][6] = 32'h45386000;
        data[46][7] = 32'h45387000;
        data[46][8] = 32'h45388000;
        data[46][9] = 32'h45389000;
        data[46][10] = 32'h4538a000;
        data[46][11] = 32'h4538b000;
        data[46][12] = 32'h4538c000;
        data[46][13] = 32'h4538d000;
        data[46][14] = 32'h4538e000;
        data[46][15] = 32'h4538f000;
        data[46][16] = 32'h45390000;
        data[46][17] = 32'h45391000;
        data[46][18] = 32'h45392000;
        data[46][19] = 32'h45393000;
        data[46][20] = 32'h45394000;
        data[46][21] = 32'h45395000;
        data[46][22] = 32'h45396000;
        data[46][23] = 32'h45397000;
        data[46][24] = 32'h45398000;
        data[46][25] = 32'h45399000;
        data[46][26] = 32'h4539a000;
        data[46][27] = 32'h4539b000;
        data[46][28] = 32'h4539c000;
        data[46][29] = 32'h4539d000;
        data[46][30] = 32'h4539e000;
        data[46][31] = 32'h4539f000;
        data[46][32] = 32'h453a0000;
        data[46][33] = 32'h453a1000;
        data[46][34] = 32'h453a2000;
        data[46][35] = 32'h453a3000;
        data[46][36] = 32'h453a4000;
        data[46][37] = 32'h453a5000;
        data[46][38] = 32'h453a6000;
        data[46][39] = 32'h453a7000;
        data[46][40] = 32'h453a8000;
        data[46][41] = 32'h453a9000;
        data[46][42] = 32'h453aa000;
        data[46][43] = 32'h453ab000;
        data[46][44] = 32'h453ac000;
        data[46][45] = 32'h453ad000;
        data[46][46] = 32'h453ae000;
        data[46][47] = 32'h453af000;
        data[46][48] = 32'h453b0000;
        data[46][49] = 32'h453b1000;
        data[46][50] = 32'h453b2000;
        data[46][51] = 32'h453b3000;
        data[46][52] = 32'h453b4000;
        data[46][53] = 32'h453b5000;
        data[46][54] = 32'h453b6000;
        data[46][55] = 32'h453b7000;
        data[46][56] = 32'h453b8000;
        data[46][57] = 32'h453b9000;
        data[46][58] = 32'h453ba000;
        data[46][59] = 32'h453bb000;
        data[46][60] = 32'h453bc000;
        data[46][61] = 32'h453bd000;
        data[46][62] = 32'h453be000;
        data[46][63] = 32'h453bf000;
        data[47][0] = 32'h453c0000;
        data[47][1] = 32'h453c1000;
        data[47][2] = 32'h453c2000;
        data[47][3] = 32'h453c3000;
        data[47][4] = 32'h453c4000;
        data[47][5] = 32'h453c5000;
        data[47][6] = 32'h453c6000;
        data[47][7] = 32'h453c7000;
        data[47][8] = 32'h453c8000;
        data[47][9] = 32'h453c9000;
        data[47][10] = 32'h453ca000;
        data[47][11] = 32'h453cb000;
        data[47][12] = 32'h453cc000;
        data[47][13] = 32'h453cd000;
        data[47][14] = 32'h453ce000;
        data[47][15] = 32'h453cf000;
        data[47][16] = 32'h453d0000;
        data[47][17] = 32'h453d1000;
        data[47][18] = 32'h453d2000;
        data[47][19] = 32'h453d3000;
        data[47][20] = 32'h453d4000;
        data[47][21] = 32'h453d5000;
        data[47][22] = 32'h453d6000;
        data[47][23] = 32'h453d7000;
        data[47][24] = 32'h453d8000;
        data[47][25] = 32'h453d9000;
        data[47][26] = 32'h453da000;
        data[47][27] = 32'h453db000;
        data[47][28] = 32'h453dc000;
        data[47][29] = 32'h453dd000;
        data[47][30] = 32'h453de000;
        data[47][31] = 32'h453df000;
        data[47][32] = 32'h453e0000;
        data[47][33] = 32'h453e1000;
        data[47][34] = 32'h453e2000;
        data[47][35] = 32'h453e3000;
        data[47][36] = 32'h453e4000;
        data[47][37] = 32'h453e5000;
        data[47][38] = 32'h453e6000;
        data[47][39] = 32'h453e7000;
        data[47][40] = 32'h453e8000;
        data[47][41] = 32'h453e9000;
        data[47][42] = 32'h453ea000;
        data[47][43] = 32'h453eb000;
        data[47][44] = 32'h453ec000;
        data[47][45] = 32'h453ed000;
        data[47][46] = 32'h453ee000;
        data[47][47] = 32'h453ef000;
        data[47][48] = 32'h453f0000;
        data[47][49] = 32'h453f1000;
        data[47][50] = 32'h453f2000;
        data[47][51] = 32'h453f3000;
        data[47][52] = 32'h453f4000;
        data[47][53] = 32'h453f5000;
        data[47][54] = 32'h453f6000;
        data[47][55] = 32'h453f7000;
        data[47][56] = 32'h453f8000;
        data[47][57] = 32'h453f9000;
        data[47][58] = 32'h453fa000;
        data[47][59] = 32'h453fb000;
        data[47][60] = 32'h453fc000;
        data[47][61] = 32'h453fd000;
        data[47][62] = 32'h453fe000;
        data[47][63] = 32'h453ff000;
        data[48][0] = 32'h45400000;
        data[48][1] = 32'h45401000;
        data[48][2] = 32'h45402000;
        data[48][3] = 32'h45403000;
        data[48][4] = 32'h45404000;
        data[48][5] = 32'h45405000;
        data[48][6] = 32'h45406000;
        data[48][7] = 32'h45407000;
        data[48][8] = 32'h45408000;
        data[48][9] = 32'h45409000;
        data[48][10] = 32'h4540a000;
        data[48][11] = 32'h4540b000;
        data[48][12] = 32'h4540c000;
        data[48][13] = 32'h4540d000;
        data[48][14] = 32'h4540e000;
        data[48][15] = 32'h4540f000;
        data[48][16] = 32'h45410000;
        data[48][17] = 32'h45411000;
        data[48][18] = 32'h45412000;
        data[48][19] = 32'h45413000;
        data[48][20] = 32'h45414000;
        data[48][21] = 32'h45415000;
        data[48][22] = 32'h45416000;
        data[48][23] = 32'h45417000;
        data[48][24] = 32'h45418000;
        data[48][25] = 32'h45419000;
        data[48][26] = 32'h4541a000;
        data[48][27] = 32'h4541b000;
        data[48][28] = 32'h4541c000;
        data[48][29] = 32'h4541d000;
        data[48][30] = 32'h4541e000;
        data[48][31] = 32'h4541f000;
        data[48][32] = 32'h45420000;
        data[48][33] = 32'h45421000;
        data[48][34] = 32'h45422000;
        data[48][35] = 32'h45423000;
        data[48][36] = 32'h45424000;
        data[48][37] = 32'h45425000;
        data[48][38] = 32'h45426000;
        data[48][39] = 32'h45427000;
        data[48][40] = 32'h45428000;
        data[48][41] = 32'h45429000;
        data[48][42] = 32'h4542a000;
        data[48][43] = 32'h4542b000;
        data[48][44] = 32'h4542c000;
        data[48][45] = 32'h4542d000;
        data[48][46] = 32'h4542e000;
        data[48][47] = 32'h4542f000;
        data[48][48] = 32'h45430000;
        data[48][49] = 32'h45431000;
        data[48][50] = 32'h45432000;
        data[48][51] = 32'h45433000;
        data[48][52] = 32'h45434000;
        data[48][53] = 32'h45435000;
        data[48][54] = 32'h45436000;
        data[48][55] = 32'h45437000;
        data[48][56] = 32'h45438000;
        data[48][57] = 32'h45439000;
        data[48][58] = 32'h4543a000;
        data[48][59] = 32'h4543b000;
        data[48][60] = 32'h4543c000;
        data[48][61] = 32'h4543d000;
        data[48][62] = 32'h4543e000;
        data[48][63] = 32'h4543f000;
        data[49][0] = 32'h45440000;
        data[49][1] = 32'h45441000;
        data[49][2] = 32'h45442000;
        data[49][3] = 32'h45443000;
        data[49][4] = 32'h45444000;
        data[49][5] = 32'h45445000;
        data[49][6] = 32'h45446000;
        data[49][7] = 32'h45447000;
        data[49][8] = 32'h45448000;
        data[49][9] = 32'h45449000;
        data[49][10] = 32'h4544a000;
        data[49][11] = 32'h4544b000;
        data[49][12] = 32'h4544c000;
        data[49][13] = 32'h4544d000;
        data[49][14] = 32'h4544e000;
        data[49][15] = 32'h4544f000;
        data[49][16] = 32'h45450000;
        data[49][17] = 32'h45451000;
        data[49][18] = 32'h45452000;
        data[49][19] = 32'h45453000;
        data[49][20] = 32'h45454000;
        data[49][21] = 32'h45455000;
        data[49][22] = 32'h45456000;
        data[49][23] = 32'h45457000;
        data[49][24] = 32'h45458000;
        data[49][25] = 32'h45459000;
        data[49][26] = 32'h4545a000;
        data[49][27] = 32'h4545b000;
        data[49][28] = 32'h4545c000;
        data[49][29] = 32'h4545d000;
        data[49][30] = 32'h4545e000;
        data[49][31] = 32'h4545f000;
        data[49][32] = 32'h45460000;
        data[49][33] = 32'h45461000;
        data[49][34] = 32'h45462000;
        data[49][35] = 32'h45463000;
        data[49][36] = 32'h45464000;
        data[49][37] = 32'h45465000;
        data[49][38] = 32'h45466000;
        data[49][39] = 32'h45467000;
        data[49][40] = 32'h45468000;
        data[49][41] = 32'h45469000;
        data[49][42] = 32'h4546a000;
        data[49][43] = 32'h4546b000;
        data[49][44] = 32'h4546c000;
        data[49][45] = 32'h4546d000;
        data[49][46] = 32'h4546e000;
        data[49][47] = 32'h4546f000;
        data[49][48] = 32'h45470000;
        data[49][49] = 32'h45471000;
        data[49][50] = 32'h45472000;
        data[49][51] = 32'h45473000;
        data[49][52] = 32'h45474000;
        data[49][53] = 32'h45475000;
        data[49][54] = 32'h45476000;
        data[49][55] = 32'h45477000;
        data[49][56] = 32'h45478000;
        data[49][57] = 32'h45479000;
        data[49][58] = 32'h4547a000;
        data[49][59] = 32'h4547b000;
        data[49][60] = 32'h4547c000;
        data[49][61] = 32'h4547d000;
        data[49][62] = 32'h4547e000;
        data[49][63] = 32'h4547f000;
        data[50][0] = 32'h45480000;
        data[50][1] = 32'h45481000;
        data[50][2] = 32'h45482000;
        data[50][3] = 32'h45483000;
        data[50][4] = 32'h45484000;
        data[50][5] = 32'h45485000;
        data[50][6] = 32'h45486000;
        data[50][7] = 32'h45487000;
        data[50][8] = 32'h45488000;
        data[50][9] = 32'h45489000;
        data[50][10] = 32'h4548a000;
        data[50][11] = 32'h4548b000;
        data[50][12] = 32'h4548c000;
        data[50][13] = 32'h4548d000;
        data[50][14] = 32'h4548e000;
        data[50][15] = 32'h4548f000;
        data[50][16] = 32'h45490000;
        data[50][17] = 32'h45491000;
        data[50][18] = 32'h45492000;
        data[50][19] = 32'h45493000;
        data[50][20] = 32'h45494000;
        data[50][21] = 32'h45495000;
        data[50][22] = 32'h45496000;
        data[50][23] = 32'h45497000;
        data[50][24] = 32'h45498000;
        data[50][25] = 32'h45499000;
        data[50][26] = 32'h4549a000;
        data[50][27] = 32'h4549b000;
        data[50][28] = 32'h4549c000;
        data[50][29] = 32'h4549d000;
        data[50][30] = 32'h4549e000;
        data[50][31] = 32'h4549f000;
        data[50][32] = 32'h454a0000;
        data[50][33] = 32'h454a1000;
        data[50][34] = 32'h454a2000;
        data[50][35] = 32'h454a3000;
        data[50][36] = 32'h454a4000;
        data[50][37] = 32'h454a5000;
        data[50][38] = 32'h454a6000;
        data[50][39] = 32'h454a7000;
        data[50][40] = 32'h454a8000;
        data[50][41] = 32'h454a9000;
        data[50][42] = 32'h454aa000;
        data[50][43] = 32'h454ab000;
        data[50][44] = 32'h454ac000;
        data[50][45] = 32'h454ad000;
        data[50][46] = 32'h454ae000;
        data[50][47] = 32'h454af000;
        data[50][48] = 32'h454b0000;
        data[50][49] = 32'h454b1000;
        data[50][50] = 32'h454b2000;
        data[50][51] = 32'h454b3000;
        data[50][52] = 32'h454b4000;
        data[50][53] = 32'h454b5000;
        data[50][54] = 32'h454b6000;
        data[50][55] = 32'h454b7000;
        data[50][56] = 32'h454b8000;
        data[50][57] = 32'h454b9000;
        data[50][58] = 32'h454ba000;
        data[50][59] = 32'h454bb000;
        data[50][60] = 32'h454bc000;
        data[50][61] = 32'h454bd000;
        data[50][62] = 32'h454be000;
        data[50][63] = 32'h454bf000;
        data[51][0] = 32'h454c0000;
        data[51][1] = 32'h454c1000;
        data[51][2] = 32'h454c2000;
        data[51][3] = 32'h454c3000;
        data[51][4] = 32'h454c4000;
        data[51][5] = 32'h454c5000;
        data[51][6] = 32'h454c6000;
        data[51][7] = 32'h454c7000;
        data[51][8] = 32'h454c8000;
        data[51][9] = 32'h454c9000;
        data[51][10] = 32'h454ca000;
        data[51][11] = 32'h454cb000;
        data[51][12] = 32'h454cc000;
        data[51][13] = 32'h454cd000;
        data[51][14] = 32'h454ce000;
        data[51][15] = 32'h454cf000;
        data[51][16] = 32'h454d0000;
        data[51][17] = 32'h454d1000;
        data[51][18] = 32'h454d2000;
        data[51][19] = 32'h454d3000;
        data[51][20] = 32'h454d4000;
        data[51][21] = 32'h454d5000;
        data[51][22] = 32'h454d6000;
        data[51][23] = 32'h454d7000;
        data[51][24] = 32'h454d8000;
        data[51][25] = 32'h454d9000;
        data[51][26] = 32'h454da000;
        data[51][27] = 32'h454db000;
        data[51][28] = 32'h454dc000;
        data[51][29] = 32'h454dd000;
        data[51][30] = 32'h454de000;
        data[51][31] = 32'h454df000;
        data[51][32] = 32'h454e0000;
        data[51][33] = 32'h454e1000;
        data[51][34] = 32'h454e2000;
        data[51][35] = 32'h454e3000;
        data[51][36] = 32'h454e4000;
        data[51][37] = 32'h454e5000;
        data[51][38] = 32'h454e6000;
        data[51][39] = 32'h454e7000;
        data[51][40] = 32'h454e8000;
        data[51][41] = 32'h454e9000;
        data[51][42] = 32'h454ea000;
        data[51][43] = 32'h454eb000;
        data[51][44] = 32'h454ec000;
        data[51][45] = 32'h454ed000;
        data[51][46] = 32'h454ee000;
        data[51][47] = 32'h454ef000;
        data[51][48] = 32'h454f0000;
        data[51][49] = 32'h454f1000;
        data[51][50] = 32'h454f2000;
        data[51][51] = 32'h454f3000;
        data[51][52] = 32'h454f4000;
        data[51][53] = 32'h454f5000;
        data[51][54] = 32'h454f6000;
        data[51][55] = 32'h454f7000;
        data[51][56] = 32'h454f8000;
        data[51][57] = 32'h454f9000;
        data[51][58] = 32'h454fa000;
        data[51][59] = 32'h454fb000;
        data[51][60] = 32'h454fc000;
        data[51][61] = 32'h454fd000;
        data[51][62] = 32'h454fe000;
        data[51][63] = 32'h454ff000;
        data[52][0] = 32'h45500000;
        data[52][1] = 32'h45501000;
        data[52][2] = 32'h45502000;
        data[52][3] = 32'h45503000;
        data[52][4] = 32'h45504000;
        data[52][5] = 32'h45505000;
        data[52][6] = 32'h45506000;
        data[52][7] = 32'h45507000;
        data[52][8] = 32'h45508000;
        data[52][9] = 32'h45509000;
        data[52][10] = 32'h4550a000;
        data[52][11] = 32'h4550b000;
        data[52][12] = 32'h4550c000;
        data[52][13] = 32'h4550d000;
        data[52][14] = 32'h4550e000;
        data[52][15] = 32'h4550f000;
        data[52][16] = 32'h45510000;
        data[52][17] = 32'h45511000;
        data[52][18] = 32'h45512000;
        data[52][19] = 32'h45513000;
        data[52][20] = 32'h45514000;
        data[52][21] = 32'h45515000;
        data[52][22] = 32'h45516000;
        data[52][23] = 32'h45517000;
        data[52][24] = 32'h45518000;
        data[52][25] = 32'h45519000;
        data[52][26] = 32'h4551a000;
        data[52][27] = 32'h4551b000;
        data[52][28] = 32'h4551c000;
        data[52][29] = 32'h4551d000;
        data[52][30] = 32'h4551e000;
        data[52][31] = 32'h4551f000;
        data[52][32] = 32'h45520000;
        data[52][33] = 32'h45521000;
        data[52][34] = 32'h45522000;
        data[52][35] = 32'h45523000;
        data[52][36] = 32'h45524000;
        data[52][37] = 32'h45525000;
        data[52][38] = 32'h45526000;
        data[52][39] = 32'h45527000;
        data[52][40] = 32'h45528000;
        data[52][41] = 32'h45529000;
        data[52][42] = 32'h4552a000;
        data[52][43] = 32'h4552b000;
        data[52][44] = 32'h4552c000;
        data[52][45] = 32'h4552d000;
        data[52][46] = 32'h4552e000;
        data[52][47] = 32'h4552f000;
        data[52][48] = 32'h45530000;
        data[52][49] = 32'h45531000;
        data[52][50] = 32'h45532000;
        data[52][51] = 32'h45533000;
        data[52][52] = 32'h45534000;
        data[52][53] = 32'h45535000;
        data[52][54] = 32'h45536000;
        data[52][55] = 32'h45537000;
        data[52][56] = 32'h45538000;
        data[52][57] = 32'h45539000;
        data[52][58] = 32'h4553a000;
        data[52][59] = 32'h4553b000;
        data[52][60] = 32'h4553c000;
        data[52][61] = 32'h4553d000;
        data[52][62] = 32'h4553e000;
        data[52][63] = 32'h4553f000;
        data[53][0] = 32'h45540000;
        data[53][1] = 32'h45541000;
        data[53][2] = 32'h45542000;
        data[53][3] = 32'h45543000;
        data[53][4] = 32'h45544000;
        data[53][5] = 32'h45545000;
        data[53][6] = 32'h45546000;
        data[53][7] = 32'h45547000;
        data[53][8] = 32'h45548000;
        data[53][9] = 32'h45549000;
        data[53][10] = 32'h4554a000;
        data[53][11] = 32'h4554b000;
        data[53][12] = 32'h4554c000;
        data[53][13] = 32'h4554d000;
        data[53][14] = 32'h4554e000;
        data[53][15] = 32'h4554f000;
        data[53][16] = 32'h45550000;
        data[53][17] = 32'h45551000;
        data[53][18] = 32'h45552000;
        data[53][19] = 32'h45553000;
        data[53][20] = 32'h45554000;
        data[53][21] = 32'h45555000;
        data[53][22] = 32'h45556000;
        data[53][23] = 32'h45557000;
        data[53][24] = 32'h45558000;
        data[53][25] = 32'h45559000;
        data[53][26] = 32'h4555a000;
        data[53][27] = 32'h4555b000;
        data[53][28] = 32'h4555c000;
        data[53][29] = 32'h4555d000;
        data[53][30] = 32'h4555e000;
        data[53][31] = 32'h4555f000;
        data[53][32] = 32'h45560000;
        data[53][33] = 32'h45561000;
        data[53][34] = 32'h45562000;
        data[53][35] = 32'h45563000;
        data[53][36] = 32'h45564000;
        data[53][37] = 32'h45565000;
        data[53][38] = 32'h45566000;
        data[53][39] = 32'h45567000;
        data[53][40] = 32'h45568000;
        data[53][41] = 32'h45569000;
        data[53][42] = 32'h4556a000;
        data[53][43] = 32'h4556b000;
        data[53][44] = 32'h4556c000;
        data[53][45] = 32'h4556d000;
        data[53][46] = 32'h4556e000;
        data[53][47] = 32'h4556f000;
        data[53][48] = 32'h45570000;
        data[53][49] = 32'h45571000;
        data[53][50] = 32'h45572000;
        data[53][51] = 32'h45573000;
        data[53][52] = 32'h45574000;
        data[53][53] = 32'h45575000;
        data[53][54] = 32'h45576000;
        data[53][55] = 32'h45577000;
        data[53][56] = 32'h45578000;
        data[53][57] = 32'h45579000;
        data[53][58] = 32'h4557a000;
        data[53][59] = 32'h4557b000;
        data[53][60] = 32'h4557c000;
        data[53][61] = 32'h4557d000;
        data[53][62] = 32'h4557e000;
        data[53][63] = 32'h4557f000;
        data[54][0] = 32'h45580000;
        data[54][1] = 32'h45581000;
        data[54][2] = 32'h45582000;
        data[54][3] = 32'h45583000;
        data[54][4] = 32'h45584000;
        data[54][5] = 32'h45585000;
        data[54][6] = 32'h45586000;
        data[54][7] = 32'h45587000;
        data[54][8] = 32'h45588000;
        data[54][9] = 32'h45589000;
        data[54][10] = 32'h4558a000;
        data[54][11] = 32'h4558b000;
        data[54][12] = 32'h4558c000;
        data[54][13] = 32'h4558d000;
        data[54][14] = 32'h4558e000;
        data[54][15] = 32'h4558f000;
        data[54][16] = 32'h45590000;
        data[54][17] = 32'h45591000;
        data[54][18] = 32'h45592000;
        data[54][19] = 32'h45593000;
        data[54][20] = 32'h45594000;
        data[54][21] = 32'h45595000;
        data[54][22] = 32'h45596000;
        data[54][23] = 32'h45597000;
        data[54][24] = 32'h45598000;
        data[54][25] = 32'h45599000;
        data[54][26] = 32'h4559a000;
        data[54][27] = 32'h4559b000;
        data[54][28] = 32'h4559c000;
        data[54][29] = 32'h4559d000;
        data[54][30] = 32'h4559e000;
        data[54][31] = 32'h4559f000;
        data[54][32] = 32'h455a0000;
        data[54][33] = 32'h455a1000;
        data[54][34] = 32'h455a2000;
        data[54][35] = 32'h455a3000;
        data[54][36] = 32'h455a4000;
        data[54][37] = 32'h455a5000;
        data[54][38] = 32'h455a6000;
        data[54][39] = 32'h455a7000;
        data[54][40] = 32'h455a8000;
        data[54][41] = 32'h455a9000;
        data[54][42] = 32'h455aa000;
        data[54][43] = 32'h455ab000;
        data[54][44] = 32'h455ac000;
        data[54][45] = 32'h455ad000;
        data[54][46] = 32'h455ae000;
        data[54][47] = 32'h455af000;
        data[54][48] = 32'h455b0000;
        data[54][49] = 32'h455b1000;
        data[54][50] = 32'h455b2000;
        data[54][51] = 32'h455b3000;
        data[54][52] = 32'h455b4000;
        data[54][53] = 32'h455b5000;
        data[54][54] = 32'h455b6000;
        data[54][55] = 32'h455b7000;
        data[54][56] = 32'h455b8000;
        data[54][57] = 32'h455b9000;
        data[54][58] = 32'h455ba000;
        data[54][59] = 32'h455bb000;
        data[54][60] = 32'h455bc000;
        data[54][61] = 32'h455bd000;
        data[54][62] = 32'h455be000;
        data[54][63] = 32'h455bf000;
        data[55][0] = 32'h455c0000;
        data[55][1] = 32'h455c1000;
        data[55][2] = 32'h455c2000;
        data[55][3] = 32'h455c3000;
        data[55][4] = 32'h455c4000;
        data[55][5] = 32'h455c5000;
        data[55][6] = 32'h455c6000;
        data[55][7] = 32'h455c7000;
        data[55][8] = 32'h455c8000;
        data[55][9] = 32'h455c9000;
        data[55][10] = 32'h455ca000;
        data[55][11] = 32'h455cb000;
        data[55][12] = 32'h455cc000;
        data[55][13] = 32'h455cd000;
        data[55][14] = 32'h455ce000;
        data[55][15] = 32'h455cf000;
        data[55][16] = 32'h455d0000;
        data[55][17] = 32'h455d1000;
        data[55][18] = 32'h455d2000;
        data[55][19] = 32'h455d3000;
        data[55][20] = 32'h455d4000;
        data[55][21] = 32'h455d5000;
        data[55][22] = 32'h455d6000;
        data[55][23] = 32'h455d7000;
        data[55][24] = 32'h455d8000;
        data[55][25] = 32'h455d9000;
        data[55][26] = 32'h455da000;
        data[55][27] = 32'h455db000;
        data[55][28] = 32'h455dc000;
        data[55][29] = 32'h455dd000;
        data[55][30] = 32'h455de000;
        data[55][31] = 32'h455df000;
        data[55][32] = 32'h455e0000;
        data[55][33] = 32'h455e1000;
        data[55][34] = 32'h455e2000;
        data[55][35] = 32'h455e3000;
        data[55][36] = 32'h455e4000;
        data[55][37] = 32'h455e5000;
        data[55][38] = 32'h455e6000;
        data[55][39] = 32'h455e7000;
        data[55][40] = 32'h455e8000;
        data[55][41] = 32'h455e9000;
        data[55][42] = 32'h455ea000;
        data[55][43] = 32'h455eb000;
        data[55][44] = 32'h455ec000;
        data[55][45] = 32'h455ed000;
        data[55][46] = 32'h455ee000;
        data[55][47] = 32'h455ef000;
        data[55][48] = 32'h455f0000;
        data[55][49] = 32'h455f1000;
        data[55][50] = 32'h455f2000;
        data[55][51] = 32'h455f3000;
        data[55][52] = 32'h455f4000;
        data[55][53] = 32'h455f5000;
        data[55][54] = 32'h455f6000;
        data[55][55] = 32'h455f7000;
        data[55][56] = 32'h455f8000;
        data[55][57] = 32'h455f9000;
        data[55][58] = 32'h455fa000;
        data[55][59] = 32'h455fb000;
        data[55][60] = 32'h455fc000;
        data[55][61] = 32'h455fd000;
        data[55][62] = 32'h455fe000;
        data[55][63] = 32'h455ff000;
        data[56][0] = 32'h45600000;
        data[56][1] = 32'h45601000;
        data[56][2] = 32'h45602000;
        data[56][3] = 32'h45603000;
        data[56][4] = 32'h45604000;
        data[56][5] = 32'h45605000;
        data[56][6] = 32'h45606000;
        data[56][7] = 32'h45607000;
        data[56][8] = 32'h45608000;
        data[56][9] = 32'h45609000;
        data[56][10] = 32'h4560a000;
        data[56][11] = 32'h4560b000;
        data[56][12] = 32'h4560c000;
        data[56][13] = 32'h4560d000;
        data[56][14] = 32'h4560e000;
        data[56][15] = 32'h4560f000;
        data[56][16] = 32'h45610000;
        data[56][17] = 32'h45611000;
        data[56][18] = 32'h45612000;
        data[56][19] = 32'h45613000;
        data[56][20] = 32'h45614000;
        data[56][21] = 32'h45615000;
        data[56][22] = 32'h45616000;
        data[56][23] = 32'h45617000;
        data[56][24] = 32'h45618000;
        data[56][25] = 32'h45619000;
        data[56][26] = 32'h4561a000;
        data[56][27] = 32'h4561b000;
        data[56][28] = 32'h4561c000;
        data[56][29] = 32'h4561d000;
        data[56][30] = 32'h4561e000;
        data[56][31] = 32'h4561f000;
        data[56][32] = 32'h45620000;
        data[56][33] = 32'h45621000;
        data[56][34] = 32'h45622000;
        data[56][35] = 32'h45623000;
        data[56][36] = 32'h45624000;
        data[56][37] = 32'h45625000;
        data[56][38] = 32'h45626000;
        data[56][39] = 32'h45627000;
        data[56][40] = 32'h45628000;
        data[56][41] = 32'h45629000;
        data[56][42] = 32'h4562a000;
        data[56][43] = 32'h4562b000;
        data[56][44] = 32'h4562c000;
        data[56][45] = 32'h4562d000;
        data[56][46] = 32'h4562e000;
        data[56][47] = 32'h4562f000;
        data[56][48] = 32'h45630000;
        data[56][49] = 32'h45631000;
        data[56][50] = 32'h45632000;
        data[56][51] = 32'h45633000;
        data[56][52] = 32'h45634000;
        data[56][53] = 32'h45635000;
        data[56][54] = 32'h45636000;
        data[56][55] = 32'h45637000;
        data[56][56] = 32'h45638000;
        data[56][57] = 32'h45639000;
        data[56][58] = 32'h4563a000;
        data[56][59] = 32'h4563b000;
        data[56][60] = 32'h4563c000;
        data[56][61] = 32'h4563d000;
        data[56][62] = 32'h4563e000;
        data[56][63] = 32'h4563f000;
        data[57][0] = 32'h45640000;
        data[57][1] = 32'h45641000;
        data[57][2] = 32'h45642000;
        data[57][3] = 32'h45643000;
        data[57][4] = 32'h45644000;
        data[57][5] = 32'h45645000;
        data[57][6] = 32'h45646000;
        data[57][7] = 32'h45647000;
        data[57][8] = 32'h45648000;
        data[57][9] = 32'h45649000;
        data[57][10] = 32'h4564a000;
        data[57][11] = 32'h4564b000;
        data[57][12] = 32'h4564c000;
        data[57][13] = 32'h4564d000;
        data[57][14] = 32'h4564e000;
        data[57][15] = 32'h4564f000;
        data[57][16] = 32'h45650000;
        data[57][17] = 32'h45651000;
        data[57][18] = 32'h45652000;
        data[57][19] = 32'h45653000;
        data[57][20] = 32'h45654000;
        data[57][21] = 32'h45655000;
        data[57][22] = 32'h45656000;
        data[57][23] = 32'h45657000;
        data[57][24] = 32'h45658000;
        data[57][25] = 32'h45659000;
        data[57][26] = 32'h4565a000;
        data[57][27] = 32'h4565b000;
        data[57][28] = 32'h4565c000;
        data[57][29] = 32'h4565d000;
        data[57][30] = 32'h4565e000;
        data[57][31] = 32'h4565f000;
        data[57][32] = 32'h45660000;
        data[57][33] = 32'h45661000;
        data[57][34] = 32'h45662000;
        data[57][35] = 32'h45663000;
        data[57][36] = 32'h45664000;
        data[57][37] = 32'h45665000;
        data[57][38] = 32'h45666000;
        data[57][39] = 32'h45667000;
        data[57][40] = 32'h45668000;
        data[57][41] = 32'h45669000;
        data[57][42] = 32'h4566a000;
        data[57][43] = 32'h4566b000;
        data[57][44] = 32'h4566c000;
        data[57][45] = 32'h4566d000;
        data[57][46] = 32'h4566e000;
        data[57][47] = 32'h4566f000;
        data[57][48] = 32'h45670000;
        data[57][49] = 32'h45671000;
        data[57][50] = 32'h45672000;
        data[57][51] = 32'h45673000;
        data[57][52] = 32'h45674000;
        data[57][53] = 32'h45675000;
        data[57][54] = 32'h45676000;
        data[57][55] = 32'h45677000;
        data[57][56] = 32'h45678000;
        data[57][57] = 32'h45679000;
        data[57][58] = 32'h4567a000;
        data[57][59] = 32'h4567b000;
        data[57][60] = 32'h4567c000;
        data[57][61] = 32'h4567d000;
        data[57][62] = 32'h4567e000;
        data[57][63] = 32'h4567f000;
        data[58][0] = 32'h45680000;
        data[58][1] = 32'h45681000;
        data[58][2] = 32'h45682000;
        data[58][3] = 32'h45683000;
        data[58][4] = 32'h45684000;
        data[58][5] = 32'h45685000;
        data[58][6] = 32'h45686000;
        data[58][7] = 32'h45687000;
        data[58][8] = 32'h45688000;
        data[58][9] = 32'h45689000;
        data[58][10] = 32'h4568a000;
        data[58][11] = 32'h4568b000;
        data[58][12] = 32'h4568c000;
        data[58][13] = 32'h4568d000;
        data[58][14] = 32'h4568e000;
        data[58][15] = 32'h4568f000;
        data[58][16] = 32'h45690000;
        data[58][17] = 32'h45691000;
        data[58][18] = 32'h45692000;
        data[58][19] = 32'h45693000;
        data[58][20] = 32'h45694000;
        data[58][21] = 32'h45695000;
        data[58][22] = 32'h45696000;
        data[58][23] = 32'h45697000;
        data[58][24] = 32'h45698000;
        data[58][25] = 32'h45699000;
        data[58][26] = 32'h4569a000;
        data[58][27] = 32'h4569b000;
        data[58][28] = 32'h4569c000;
        data[58][29] = 32'h4569d000;
        data[58][30] = 32'h4569e000;
        data[58][31] = 32'h4569f000;
        data[58][32] = 32'h456a0000;
        data[58][33] = 32'h456a1000;
        data[58][34] = 32'h456a2000;
        data[58][35] = 32'h456a3000;
        data[58][36] = 32'h456a4000;
        data[58][37] = 32'h456a5000;
        data[58][38] = 32'h456a6000;
        data[58][39] = 32'h456a7000;
        data[58][40] = 32'h456a8000;
        data[58][41] = 32'h456a9000;
        data[58][42] = 32'h456aa000;
        data[58][43] = 32'h456ab000;
        data[58][44] = 32'h456ac000;
        data[58][45] = 32'h456ad000;
        data[58][46] = 32'h456ae000;
        data[58][47] = 32'h456af000;
        data[58][48] = 32'h456b0000;
        data[58][49] = 32'h456b1000;
        data[58][50] = 32'h456b2000;
        data[58][51] = 32'h456b3000;
        data[58][52] = 32'h456b4000;
        data[58][53] = 32'h456b5000;
        data[58][54] = 32'h456b6000;
        data[58][55] = 32'h456b7000;
        data[58][56] = 32'h456b8000;
        data[58][57] = 32'h456b9000;
        data[58][58] = 32'h456ba000;
        data[58][59] = 32'h456bb000;
        data[58][60] = 32'h456bc000;
        data[58][61] = 32'h456bd000;
        data[58][62] = 32'h456be000;
        data[58][63] = 32'h456bf000;
        data[59][0] = 32'h456c0000;
        data[59][1] = 32'h456c1000;
        data[59][2] = 32'h456c2000;
        data[59][3] = 32'h456c3000;
        data[59][4] = 32'h456c4000;
        data[59][5] = 32'h456c5000;
        data[59][6] = 32'h456c6000;
        data[59][7] = 32'h456c7000;
        data[59][8] = 32'h456c8000;
        data[59][9] = 32'h456c9000;
        data[59][10] = 32'h456ca000;
        data[59][11] = 32'h456cb000;
        data[59][12] = 32'h456cc000;
        data[59][13] = 32'h456cd000;
        data[59][14] = 32'h456ce000;
        data[59][15] = 32'h456cf000;
        data[59][16] = 32'h456d0000;
        data[59][17] = 32'h456d1000;
        data[59][18] = 32'h456d2000;
        data[59][19] = 32'h456d3000;
        data[59][20] = 32'h456d4000;
        data[59][21] = 32'h456d5000;
        data[59][22] = 32'h456d6000;
        data[59][23] = 32'h456d7000;
        data[59][24] = 32'h456d8000;
        data[59][25] = 32'h456d9000;
        data[59][26] = 32'h456da000;
        data[59][27] = 32'h456db000;
        data[59][28] = 32'h456dc000;
        data[59][29] = 32'h456dd000;
        data[59][30] = 32'h456de000;
        data[59][31] = 32'h456df000;
        data[59][32] = 32'h456e0000;
        data[59][33] = 32'h456e1000;
        data[59][34] = 32'h456e2000;
        data[59][35] = 32'h456e3000;
        data[59][36] = 32'h456e4000;
        data[59][37] = 32'h456e5000;
        data[59][38] = 32'h456e6000;
        data[59][39] = 32'h456e7000;
        data[59][40] = 32'h456e8000;
        data[59][41] = 32'h456e9000;
        data[59][42] = 32'h456ea000;
        data[59][43] = 32'h456eb000;
        data[59][44] = 32'h456ec000;
        data[59][45] = 32'h456ed000;
        data[59][46] = 32'h456ee000;
        data[59][47] = 32'h456ef000;
        data[59][48] = 32'h456f0000;
        data[59][49] = 32'h456f1000;
        data[59][50] = 32'h456f2000;
        data[59][51] = 32'h456f3000;
        data[59][52] = 32'h456f4000;
        data[59][53] = 32'h456f5000;
        data[59][54] = 32'h456f6000;
        data[59][55] = 32'h456f7000;
        data[59][56] = 32'h456f8000;
        data[59][57] = 32'h456f9000;
        data[59][58] = 32'h456fa000;
        data[59][59] = 32'h456fb000;
        data[59][60] = 32'h456fc000;
        data[59][61] = 32'h456fd000;
        data[59][62] = 32'h456fe000;
        data[59][63] = 32'h456ff000;
        data[60][0] = 32'h45700000;
        data[60][1] = 32'h45701000;
        data[60][2] = 32'h45702000;
        data[60][3] = 32'h45703000;
        data[60][4] = 32'h45704000;
        data[60][5] = 32'h45705000;
        data[60][6] = 32'h45706000;
        data[60][7] = 32'h45707000;
        data[60][8] = 32'h45708000;
        data[60][9] = 32'h45709000;
        data[60][10] = 32'h4570a000;
        data[60][11] = 32'h4570b000;
        data[60][12] = 32'h4570c000;
        data[60][13] = 32'h4570d000;
        data[60][14] = 32'h4570e000;
        data[60][15] = 32'h4570f000;
        data[60][16] = 32'h45710000;
        data[60][17] = 32'h45711000;
        data[60][18] = 32'h45712000;
        data[60][19] = 32'h45713000;
        data[60][20] = 32'h45714000;
        data[60][21] = 32'h45715000;
        data[60][22] = 32'h45716000;
        data[60][23] = 32'h45717000;
        data[60][24] = 32'h45718000;
        data[60][25] = 32'h45719000;
        data[60][26] = 32'h4571a000;
        data[60][27] = 32'h4571b000;
        data[60][28] = 32'h4571c000;
        data[60][29] = 32'h4571d000;
        data[60][30] = 32'h4571e000;
        data[60][31] = 32'h4571f000;
        data[60][32] = 32'h45720000;
        data[60][33] = 32'h45721000;
        data[60][34] = 32'h45722000;
        data[60][35] = 32'h45723000;
        data[60][36] = 32'h45724000;
        data[60][37] = 32'h45725000;
        data[60][38] = 32'h45726000;
        data[60][39] = 32'h45727000;
        data[60][40] = 32'h45728000;
        data[60][41] = 32'h45729000;
        data[60][42] = 32'h4572a000;
        data[60][43] = 32'h4572b000;
        data[60][44] = 32'h4572c000;
        data[60][45] = 32'h4572d000;
        data[60][46] = 32'h4572e000;
        data[60][47] = 32'h4572f000;
        data[60][48] = 32'h45730000;
        data[60][49] = 32'h45731000;
        data[60][50] = 32'h45732000;
        data[60][51] = 32'h45733000;
        data[60][52] = 32'h45734000;
        data[60][53] = 32'h45735000;
        data[60][54] = 32'h45736000;
        data[60][55] = 32'h45737000;
        data[60][56] = 32'h45738000;
        data[60][57] = 32'h45739000;
        data[60][58] = 32'h4573a000;
        data[60][59] = 32'h4573b000;
        data[60][60] = 32'h4573c000;
        data[60][61] = 32'h4573d000;
        data[60][62] = 32'h4573e000;
        data[60][63] = 32'h4573f000;
        data[61][0] = 32'h45740000;
        data[61][1] = 32'h45741000;
        data[61][2] = 32'h45742000;
        data[61][3] = 32'h45743000;
        data[61][4] = 32'h45744000;
        data[61][5] = 32'h45745000;
        data[61][6] = 32'h45746000;
        data[61][7] = 32'h45747000;
        data[61][8] = 32'h45748000;
        data[61][9] = 32'h45749000;
        data[61][10] = 32'h4574a000;
        data[61][11] = 32'h4574b000;
        data[61][12] = 32'h4574c000;
        data[61][13] = 32'h4574d000;
        data[61][14] = 32'h4574e000;
        data[61][15] = 32'h4574f000;
        data[61][16] = 32'h45750000;
        data[61][17] = 32'h45751000;
        data[61][18] = 32'h45752000;
        data[61][19] = 32'h45753000;
        data[61][20] = 32'h45754000;
        data[61][21] = 32'h45755000;
        data[61][22] = 32'h45756000;
        data[61][23] = 32'h45757000;
        data[61][24] = 32'h45758000;
        data[61][25] = 32'h45759000;
        data[61][26] = 32'h4575a000;
        data[61][27] = 32'h4575b000;
        data[61][28] = 32'h4575c000;
        data[61][29] = 32'h4575d000;
        data[61][30] = 32'h4575e000;
        data[61][31] = 32'h4575f000;
        data[61][32] = 32'h45760000;
        data[61][33] = 32'h45761000;
        data[61][34] = 32'h45762000;
        data[61][35] = 32'h45763000;
        data[61][36] = 32'h45764000;
        data[61][37] = 32'h45765000;
        data[61][38] = 32'h45766000;
        data[61][39] = 32'h45767000;
        data[61][40] = 32'h45768000;
        data[61][41] = 32'h45769000;
        data[61][42] = 32'h4576a000;
        data[61][43] = 32'h4576b000;
        data[61][44] = 32'h4576c000;
        data[61][45] = 32'h4576d000;
        data[61][46] = 32'h4576e000;
        data[61][47] = 32'h4576f000;
        data[61][48] = 32'h45770000;
        data[61][49] = 32'h45771000;
        data[61][50] = 32'h45772000;
        data[61][51] = 32'h45773000;
        data[61][52] = 32'h45774000;
        data[61][53] = 32'h45775000;
        data[61][54] = 32'h45776000;
        data[61][55] = 32'h45777000;
        data[61][56] = 32'h45778000;
        data[61][57] = 32'h45779000;
        data[61][58] = 32'h4577a000;
        data[61][59] = 32'h4577b000;
        data[61][60] = 32'h4577c000;
        data[61][61] = 32'h4577d000;
        data[61][62] = 32'h4577e000;
        data[61][63] = 32'h4577f000;
        data[62][0] = 32'h45780000;
        data[62][1] = 32'h45781000;
        data[62][2] = 32'h45782000;
        data[62][3] = 32'h45783000;
        data[62][4] = 32'h45784000;
        data[62][5] = 32'h45785000;
        data[62][6] = 32'h45786000;
        data[62][7] = 32'h45787000;
        data[62][8] = 32'h45788000;
        data[62][9] = 32'h45789000;
        data[62][10] = 32'h4578a000;
        data[62][11] = 32'h4578b000;
        data[62][12] = 32'h4578c000;
        data[62][13] = 32'h4578d000;
        data[62][14] = 32'h4578e000;
        data[62][15] = 32'h4578f000;
        data[62][16] = 32'h45790000;
        data[62][17] = 32'h45791000;
        data[62][18] = 32'h45792000;
        data[62][19] = 32'h45793000;
        data[62][20] = 32'h45794000;
        data[62][21] = 32'h45795000;
        data[62][22] = 32'h45796000;
        data[62][23] = 32'h45797000;
        data[62][24] = 32'h45798000;
        data[62][25] = 32'h45799000;
        data[62][26] = 32'h4579a000;
        data[62][27] = 32'h4579b000;
        data[62][28] = 32'h4579c000;
        data[62][29] = 32'h4579d000;
        data[62][30] = 32'h4579e000;
        data[62][31] = 32'h4579f000;
        data[62][32] = 32'h457a0000;
        data[62][33] = 32'h457a1000;
        data[62][34] = 32'h457a2000;
        data[62][35] = 32'h457a3000;
        data[62][36] = 32'h457a4000;
        data[62][37] = 32'h457a5000;
        data[62][38] = 32'h457a6000;
        data[62][39] = 32'h457a7000;
        data[62][40] = 32'h457a8000;
        data[62][41] = 32'h457a9000;
        data[62][42] = 32'h457aa000;
        data[62][43] = 32'h457ab000;
        data[62][44] = 32'h457ac000;
        data[62][45] = 32'h457ad000;
        data[62][46] = 32'h457ae000;
        data[62][47] = 32'h457af000;
        data[62][48] = 32'h457b0000;
        data[62][49] = 32'h457b1000;
        data[62][50] = 32'h457b2000;
        data[62][51] = 32'h457b3000;
        data[62][52] = 32'h457b4000;
        data[62][53] = 32'h457b5000;
        data[62][54] = 32'h457b6000;
        data[62][55] = 32'h457b7000;
        data[62][56] = 32'h457b8000;
        data[62][57] = 32'h457b9000;
        data[62][58] = 32'h457ba000;
        data[62][59] = 32'h457bb000;
        data[62][60] = 32'h457bc000;
        data[62][61] = 32'h457bd000;
        data[62][62] = 32'h457be000;
        data[62][63] = 32'h457bf000;
        data[63][0] = 32'h457c0000;
        data[63][1] = 32'h457c1000;
        data[63][2] = 32'h457c2000;
        data[63][3] = 32'h457c3000;
        data[63][4] = 32'h457c4000;
        data[63][5] = 32'h457c5000;
        data[63][6] = 32'h457c6000;
        data[63][7] = 32'h457c7000;
        data[63][8] = 32'h457c8000;
        data[63][9] = 32'h457c9000;
        data[63][10] = 32'h457ca000;
        data[63][11] = 32'h457cb000;
        data[63][12] = 32'h457cc000;
        data[63][13] = 32'h457cd000;
        data[63][14] = 32'h457ce000;
        data[63][15] = 32'h457cf000;
        data[63][16] = 32'h457d0000;
        data[63][17] = 32'h457d1000;
        data[63][18] = 32'h457d2000;
        data[63][19] = 32'h457d3000;
        data[63][20] = 32'h457d4000;
        data[63][21] = 32'h457d5000;
        data[63][22] = 32'h457d6000;
        data[63][23] = 32'h457d7000;
        data[63][24] = 32'h457d8000;
        data[63][25] = 32'h457d9000;
        data[63][26] = 32'h457da000;
        data[63][27] = 32'h457db000;
        data[63][28] = 32'h457dc000;
        data[63][29] = 32'h457dd000;
        data[63][30] = 32'h457de000;
        data[63][31] = 32'h457df000;
        data[63][32] = 32'h457e0000;
        data[63][33] = 32'h457e1000;
        data[63][34] = 32'h457e2000;
        data[63][35] = 32'h457e3000;
        data[63][36] = 32'h457e4000;
        data[63][37] = 32'h457e5000;
        data[63][38] = 32'h457e6000;
        data[63][39] = 32'h457e7000;
        data[63][40] = 32'h457e8000;
        data[63][41] = 32'h457e9000;
        data[63][42] = 32'h457ea000;
        data[63][43] = 32'h457eb000;
        data[63][44] = 32'h457ec000;
        data[63][45] = 32'h457ed000;
        data[63][46] = 32'h457ee000;
        data[63][47] = 32'h457ef000;
        data[63][48] = 32'h457f0000;
        data[63][49] = 32'h457f1000;
        data[63][50] = 32'h457f2000;
        data[63][51] = 32'h457f3000;
        data[63][52] = 32'h457f4000;
        data[63][53] = 32'h457f5000;
        data[63][54] = 32'h457f6000;
        data[63][55] = 32'h457f7000;
        data[63][56] = 32'h457f8000;
        data[63][57] = 32'h457f9000;
        data[63][58] = 32'h457fa000;
        data[63][59] = 32'h457fb000;
        data[63][60] = 32'h457fc000;
        data[63][61] = 32'h457fd000;
        data[63][62] = 32'h457fe000;
        data[63][63] = 32'h457ff000;
	end
	
	
	
	// Assign output
	always @(posedge clk) begin
		if (reset) begin
			for (int i = 0; i < 64; i++) begin
				row_reg[i] <= 32'h00000000;
         end
		end else begin
			for (int i = 0; i < 4; i++) begin
				row_reg[i]    <= data[row_sel][0  + i * 16];
				row_reg[i+4]  <= data[row_sel][4  + i * 16];
				row_reg[i+8]  <= data[row_sel][8  + i * 16];
				row_reg[i+12] <= data[row_sel][12 + i * 16];
				
				row_reg[i+16] <= data[row_sel][1  + i * 16];
				row_reg[i+20] <= data[row_sel][5  + i * 16];
				row_reg[i+24] <= data[row_sel][9  + i * 16];
				row_reg[i+28] <= data[row_sel][13 + i * 16];
				
				row_reg[i+32] <= data[row_sel][2  + i * 16];
				row_reg[i+36] <= data[row_sel][6  + i * 16];
				row_reg[i+40] <= data[row_sel][10 + i * 16];
				row_reg[i+44] <= data[row_sel][14 + i * 16];
				
				row_reg[i+48] <= data[row_sel][3  + i * 16];
				row_reg[i+52] <= data[row_sel][7  + i * 16];
				row_reg[i+56] <= data[row_sel][11 + i * 16];
				row_reg[i+60] <= data[row_sel][15 + i * 16];
			end
		end
	end
	assign row = row_reg;

endmodule
