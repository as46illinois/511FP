module w64_rom
(
	output logic[31:0] w64r[63:0],
	output logic[31:0] w64i[63:0]
);

	initial begin
		w64r[0] = 32'h3f800000;
		w64i[0] = 32'h00000000;
		w64r[1] = 32'h3f800000;
		w64i[1] = 32'h00000000;
		w64r[2] = 32'h3f800000;
		w64i[2] = 32'h00000000;
		w64r[3] = 32'h3f800000;
		w64i[3] = 32'h00000000;
		w64r[4] = 32'h3f800000;
		w64i[4] = 32'h00000000;
		w64r[5] = 32'h3f800000;
		w64i[5] = 32'h00000000;
		w64r[6] = 32'h3f800000;
		w64i[6] = 32'h00000000;
		w64r[7] = 32'h3f800000;
		w64i[7] = 32'h00000000;
		w64r[8] = 32'h3f800000;
		w64i[8] = 32'h00000000;
		w64r[9] = 32'h3f800000;
		w64i[9] = 32'h00000000;
		w64r[10] = 32'h3f800000;
		w64i[10] = 32'h00000000;
		w64r[11] = 32'h3f800000;
		w64i[11] = 32'h00000000;
		w64r[12] = 32'h3f800000;
		w64i[12] = 32'h00000000;
		w64r[13] = 32'h3f800000;
		w64i[13] = 32'h00000000;
		w64r[14] = 32'h3f800000;
		w64i[14] = 32'h00000000;
		w64r[15] = 32'h3f800000;
		w64i[15] = 32'h00000000;
		w64r[16] = 32'h3f800000;
		w64i[16] = 32'h00000000;
		w64r[17] = 32'h3f7ec46d;
		w64i[17] = 32'hbdc8bd36;
		w64r[18] = 32'h3f7b14be;
		w64i[18] = 32'hbe47c5c2;
		w64r[19] = 32'h3f74fa0b;
		w64i[19] = 32'hbe94a031;
		w64r[20] = 32'h3f6c835e;
		w64i[20] = 32'hbec3ef15;
		w64r[21] = 32'h3f61c598;
		w64i[21] = 32'hbef15aea;
		w64r[22] = 32'h3f54db31;
		w64i[22] = 32'hbf0e39da;
		w64r[23] = 32'h3f45e403;
		w64i[23] = 32'hbf226799;
		w64r[24] = 32'h3f3504f3;
		w64i[24] = 32'hbf3504f3;
		w64r[25] = 32'h3f226799;
		w64i[25] = 32'hbf45e403;
		w64r[26] = 32'h3f0e39da;
		w64i[26] = 32'hbf54db31;
		w64r[27] = 32'h3ef15aea;
		w64i[27] = 32'hbf61c598;
		w64r[28] = 32'h3ec3ef15;
		w64i[28] = 32'hbf6c835e;
		w64r[29] = 32'h3e94a031;
		w64i[29] = 32'hbf74fa0b;
		w64r[30] = 32'h3e47c5c2;
		w64i[30] = 32'hbf7b14be;
		w64r[31] = 32'h3dc8bd36;
		w64i[31] = 32'hbf7ec46d;
		w64r[32] = 32'h3f800000;
		w64i[32] = 32'h00000000;
		w64r[33] = 32'h3f7b14be;
		w64i[33] = 32'hbe47c5c2;
		w64r[34] = 32'h3f6c835e;
		w64i[34] = 32'hbec3ef15;
		w64r[35] = 32'h3f54db31;
		w64i[35] = 32'hbf0e39da;
		w64r[36] = 32'h3f3504f3;
		w64i[36] = 32'hbf3504f3;
		w64r[37] = 32'h3f0e39da;
		w64i[37] = 32'hbf54db31;
		w64r[38] = 32'h3ec3ef15;
		w64i[38] = 32'hbf6c835e;
		w64r[39] = 32'h3e47c5c2;
		w64i[39] = 32'hbf7b14be;
		w64r[40] = 32'h248d3132;
		w64i[40] = 32'hbf800000;
		w64r[41] = 32'hbe47c5c2;
		w64i[41] = 32'hbf7b14be;
		w64r[42] = 32'hbec3ef15;
		w64i[42] = 32'hbf6c835e;
		w64r[43] = 32'hbf0e39da;
		w64i[43] = 32'hbf54db31;
		w64r[44] = 32'hbf3504f3;
		w64i[44] = 32'hbf3504f3;
		w64r[45] = 32'hbf54db31;
		w64i[45] = 32'hbf0e39da;
		w64r[46] = 32'hbf6c835e;
		w64i[46] = 32'hbec3ef15;
		w64r[47] = 32'hbf7b14be;
		w64i[47] = 32'hbe47c5c2;
		w64r[48] = 32'h3f800000;
		w64i[48] = 32'h00000000;
		w64r[49] = 32'h3f74fa0b;
		w64i[49] = 32'hbe94a031;
		w64r[50] = 32'h3f54db31;
		w64i[50] = 32'hbf0e39da;
		w64r[51] = 32'h3f226799;
		w64i[51] = 32'hbf45e403;
		w64r[52] = 32'h3ec3ef15;
		w64i[52] = 32'hbf6c835e;
		w64r[53] = 32'h3dc8bd36;
		w64i[53] = 32'hbf7ec46d;
		w64r[54] = 32'hbe47c5c2;
		w64i[54] = 32'hbf7b14be;
		w64r[55] = 32'hbef15aea;
		w64i[55] = 32'hbf61c598;
		w64r[56] = 32'hbf3504f3;
		w64i[56] = 32'hbf3504f3;
		w64r[57] = 32'hbf61c598;
		w64i[57] = 32'hbef15aea;
		w64r[58] = 32'hbf7b14be;
		w64i[58] = 32'hbe47c5c2;
		w64r[59] = 32'hbf7ec46d;
		w64i[59] = 32'h3dc8bd36;
		w64r[60] = 32'hbf6c835e;
		w64i[60] = 32'h3ec3ef15;
		w64r[61] = 32'hbf45e403;
		w64i[61] = 32'h3f226799;
		w64r[62] = 32'hbf0e39da;
		w64i[62] = 32'h3f54db31;
		w64r[63] = 32'hbe94a031;
		w64i[63] = 32'h3f74fa0b;
	end

endmodule
